magic
tech sky130A
magscale 1 2
timestamp 1686145127
<< obsli1 >>
rect 1104 2159 58880 57681
<< obsm1 >>
rect 934 2128 58958 57712
<< metal2 >>
rect 938 59200 994 60000
rect 2870 59200 2926 60000
rect 4802 59200 4858 60000
rect 6734 59200 6790 60000
rect 8666 59200 8722 60000
rect 10598 59200 10654 60000
rect 12530 59200 12586 60000
rect 14462 59200 14518 60000
rect 16394 59200 16450 60000
rect 18326 59200 18382 60000
rect 20258 59200 20314 60000
rect 22190 59200 22246 60000
rect 24122 59200 24178 60000
rect 26054 59200 26110 60000
rect 27986 59200 28042 60000
rect 29918 59200 29974 60000
rect 31850 59200 31906 60000
rect 33782 59200 33838 60000
rect 35714 59200 35770 60000
rect 37646 59200 37702 60000
rect 39578 59200 39634 60000
rect 41510 59200 41566 60000
rect 43442 59200 43498 60000
rect 45374 59200 45430 60000
rect 47306 59200 47362 60000
rect 49238 59200 49294 60000
rect 51170 59200 51226 60000
rect 53102 59200 53158 60000
rect 55034 59200 55090 60000
rect 56966 59200 57022 60000
rect 58898 59200 58954 60000
<< obsm2 >>
rect 1050 59144 2814 59242
rect 2982 59144 4746 59242
rect 4914 59144 6678 59242
rect 6846 59144 8610 59242
rect 8778 59144 10542 59242
rect 10710 59144 12474 59242
rect 12642 59144 14406 59242
rect 14574 59144 16338 59242
rect 16506 59144 18270 59242
rect 18438 59144 20202 59242
rect 20370 59144 22134 59242
rect 22302 59144 24066 59242
rect 24234 59144 25998 59242
rect 26166 59144 27930 59242
rect 28098 59144 29862 59242
rect 30030 59144 31794 59242
rect 31962 59144 33726 59242
rect 33894 59144 35658 59242
rect 35826 59144 37590 59242
rect 37758 59144 39522 59242
rect 39690 59144 41454 59242
rect 41622 59144 43386 59242
rect 43554 59144 45318 59242
rect 45486 59144 47250 59242
rect 47418 59144 49182 59242
rect 49350 59144 51114 59242
rect 51282 59144 53046 59242
rect 53214 59144 54978 59242
rect 55146 59144 56910 59242
rect 57078 59144 58842 59242
rect 940 2139 58952 59144
<< metal3 >>
rect 59200 44888 60000 45008
rect 59200 14968 60000 15088
<< obsm3 >>
rect 2346 45088 59200 57697
rect 2346 44808 59120 45088
rect 2346 15168 59200 44808
rect 2346 14888 59120 15168
rect 2346 2143 59200 14888
<< metal4 >>
rect 2344 2128 2664 57712
rect 3004 2128 3324 57712
rect 33064 2128 33384 57712
rect 33724 2128 34044 57712
<< metal5 >>
rect 1056 34712 58928 35032
rect 1056 34052 58928 34372
rect 1056 4076 58928 4396
rect 1056 3416 58928 3736
<< labels >>
rlabel metal5 s 1056 34712 58928 35032 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 4076 58928 4396 6 VGND
port 1 nsew ground default
rlabel metal4 s 33724 2128 34044 57712 6 VGND
port 1 nsew ground default
rlabel metal4 s 3004 2128 3324 57712 6 VGND
port 1 nsew ground default
rlabel metal5 s 1056 34052 58928 34372 6 VPWR
port 2 nsew power default
rlabel metal5 s 1056 3416 58928 3736 6 VPWR
port 2 nsew power default
rlabel metal4 s 33064 2128 33384 57712 6 VPWR
port 2 nsew power default
rlabel metal4 s 2344 2128 2664 57712 6 VPWR
port 2 nsew power default
rlabel metal3 s 59200 14968 60000 15088 6 clk
port 3 nsew
rlabel metal3 s 59200 44888 60000 45008 6 reset
port 4 nsew
rlabel metal2 s 938 59200 994 60000 6 scan_in
port 5 nsew
rlabel metal2 s 2870 59200 2926 60000 6 scan_out[0]
port 6 nsew
rlabel metal2 s 22190 59200 22246 60000 6 scan_out[10]
port 7 nsew
rlabel metal2 s 24122 59200 24178 60000 6 scan_out[11]
port 8 nsew
rlabel metal2 s 26054 59200 26110 60000 6 scan_out[12]
port 9 nsew
rlabel metal2 s 27986 59200 28042 60000 6 scan_out[13]
port 10 nsew
rlabel metal2 s 29918 59200 29974 60000 6 scan_out[14]
port 11 nsew
rlabel metal2 s 31850 59200 31906 60000 6 scan_out[15]
port 12 nsew
rlabel metal2 s 33782 59200 33838 60000 6 scan_out[16]
port 13 nsew
rlabel metal2 s 35714 59200 35770 60000 6 scan_out[17]
port 14 nsew
rlabel metal2 s 37646 59200 37702 60000 6 scan_out[18]
port 15 nsew
rlabel metal2 s 39578 59200 39634 60000 6 scan_out[19]
port 16 nsew
rlabel metal2 s 4802 59200 4858 60000 6 scan_out[1]
port 17 nsew
rlabel metal2 s 41510 59200 41566 60000 6 scan_out[20]
port 18 nsew
rlabel metal2 s 43442 59200 43498 60000 6 scan_out[21]
port 19 nsew
rlabel metal2 s 45374 59200 45430 60000 6 scan_out[22]
port 20 nsew
rlabel metal2 s 47306 59200 47362 60000 6 scan_out[23]
port 21 nsew
rlabel metal2 s 49238 59200 49294 60000 6 scan_out[24]
port 22 nsew
rlabel metal2 s 51170 59200 51226 60000 6 scan_out[25]
port 23 nsew
rlabel metal2 s 53102 59200 53158 60000 6 scan_out[26]
port 24 nsew
rlabel metal2 s 55034 59200 55090 60000 6 scan_out[27]
port 25 nsew
rlabel metal2 s 56966 59200 57022 60000 6 scan_out[28]
port 26 nsew
rlabel metal2 s 58898 59200 58954 60000 6 scan_out[29]
port 27 nsew
rlabel metal2 s 6734 59200 6790 60000 6 scan_out[2]
port 28 nsew
rlabel metal2 s 8666 59200 8722 60000 6 scan_out[3]
port 29 nsew
rlabel metal2 s 10598 59200 10654 60000 6 scan_out[4]
port 30 nsew
rlabel metal2 s 12530 59200 12586 60000 6 scan_out[5]
port 31 nsew
rlabel metal2 s 14462 59200 14518 60000 6 scan_out[6]
port 32 nsew
rlabel metal2 s 16394 59200 16450 60000 6 scan_out[7]
port 33 nsew
rlabel metal2 s 18326 59200 18382 60000 6 scan_out[8]
port 34 nsew
rlabel metal2 s 20258 59200 20314 60000 6 scan_out[9]
port 35 nsew
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1191708
string GDS_FILE /openlane/designs/scan/runs/RUN_2023.06.07_13.37.15/results/signoff/scan_chain.magic.gds
string GDS_START 87756
<< end >>

