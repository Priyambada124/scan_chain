magic
tech sky130A
magscale 1 2
timestamp 1686145206
<< checkpaint >>
rect -2998 -1804 63932 63932
<< viali >>
rect 6929 57545 6963 57579
rect 26249 57545 26283 57579
rect 28273 57545 28307 57579
rect 30389 57545 30423 57579
rect 34161 57545 34195 57579
rect 35909 57545 35943 57579
rect 45661 57545 45695 57579
rect 47777 57545 47811 57579
rect 49709 57545 49743 57579
rect 51457 57545 51491 57579
rect 53389 57545 53423 57579
rect 55505 57545 55539 57579
rect 57253 57545 57287 57579
rect 2973 57477 3007 57511
rect 4905 57477 4939 57511
rect 8953 57477 8987 57511
rect 10701 57477 10735 57511
rect 11069 57477 11103 57511
rect 12633 57477 12667 57511
rect 14565 57477 14599 57511
rect 16681 57477 16715 57511
rect 18429 57477 18463 57511
rect 20361 57477 20395 57511
rect 22293 57477 22327 57511
rect 24409 57477 24443 57511
rect 32137 57477 32171 57511
rect 37749 57477 37783 57511
rect 39865 57477 39899 57511
rect 41613 57477 41647 57511
rect 43545 57477 43579 57511
rect 55413 57477 55447 57511
rect 58173 57477 58207 57511
rect 58541 57477 58575 57511
rect 1409 57409 1443 57443
rect 3341 57409 3375 57443
rect 5273 57409 5307 57443
rect 7205 57409 7239 57443
rect 9321 57409 9355 57443
rect 13001 57409 13035 57443
rect 14933 57409 14967 57443
rect 17049 57409 17083 57443
rect 18797 57409 18831 57443
rect 20729 57409 20763 57443
rect 22661 57409 22695 57443
rect 24777 57409 24811 57443
rect 26525 57409 26559 57443
rect 28181 57409 28215 57443
rect 30113 57409 30147 57443
rect 32505 57409 32539 57443
rect 34253 57409 34287 57443
rect 36185 57409 36219 57443
rect 38117 57409 38151 57443
rect 40233 57409 40267 57443
rect 41981 57409 42015 57443
rect 43913 57409 43947 57443
rect 45569 57409 45603 57443
rect 47685 57409 47719 57443
rect 49433 57409 49467 57443
rect 51365 57409 51399 57443
rect 53297 57409 53331 57443
rect 57161 57409 57195 57443
rect 1685 57341 1719 57375
rect 16865 57001 16899 57035
rect 15853 56933 15887 56967
rect 52561 56933 52595 56967
rect 16405 56865 16439 56899
rect 17509 56865 17543 56899
rect 21925 56865 21959 56899
rect 51825 56865 51859 56899
rect 52009 56865 52043 56899
rect 53021 56865 53055 56899
rect 53113 56865 53147 56899
rect 15577 56797 15611 56831
rect 16221 56797 16255 56831
rect 16681 56797 16715 56831
rect 17785 56797 17819 56831
rect 18337 56797 18371 56831
rect 22201 56797 22235 56831
rect 23029 56797 23063 56831
rect 27077 56797 27111 56831
rect 27813 56797 27847 56831
rect 28181 56797 28215 56831
rect 51457 56797 51491 56831
rect 16313 56729 16347 56763
rect 17325 56729 17359 56763
rect 18061 56729 18095 56763
rect 52101 56729 52135 56763
rect 15761 56661 15795 56695
rect 16957 56661 16991 56695
rect 17417 56661 17451 56695
rect 18521 56661 18555 56695
rect 20453 56661 20487 56695
rect 23673 56661 23707 56695
rect 26525 56661 26559 56695
rect 27261 56661 27295 56695
rect 27997 56661 28031 56695
rect 51641 56661 51675 56695
rect 52469 56661 52503 56695
rect 52929 56661 52963 56695
rect 15209 56457 15243 56491
rect 15301 56457 15335 56491
rect 16221 56457 16255 56491
rect 17877 56457 17911 56491
rect 23489 56457 23523 56491
rect 23949 56457 23983 56491
rect 25145 56457 25179 56491
rect 26341 56457 26375 56491
rect 26801 56457 26835 56491
rect 28181 56457 28215 56491
rect 32137 56457 32171 56491
rect 32597 56457 32631 56491
rect 34713 56457 34747 56491
rect 36645 56457 36679 56491
rect 38393 56457 38427 56491
rect 38485 56457 38519 56491
rect 40325 56457 40359 56491
rect 42441 56457 42475 56491
rect 49249 56457 49283 56491
rect 49801 56457 49835 56491
rect 51457 56457 51491 56491
rect 52745 56457 52779 56491
rect 16129 56389 16163 56423
rect 16957 56389 16991 56423
rect 21373 56389 21407 56423
rect 23581 56389 23615 56423
rect 25237 56389 25271 56423
rect 27721 56389 27755 56423
rect 42809 56389 42843 56423
rect 44465 56389 44499 56423
rect 45385 56389 45419 56423
rect 49341 56389 49375 56423
rect 51365 56389 51399 56423
rect 53205 56389 53239 56423
rect 17785 56321 17819 56355
rect 18613 56321 18647 56355
rect 19441 56321 19475 56355
rect 22201 56321 22235 56355
rect 22845 56321 22879 56355
rect 24225 56321 24259 56355
rect 25881 56305 25915 56339
rect 26433 56321 26467 56355
rect 27169 56321 27203 56355
rect 27813 56321 27847 56355
rect 28641 56321 28675 56355
rect 31769 56321 31803 56355
rect 32505 56321 32539 56355
rect 34345 56321 34379 56355
rect 34989 56321 35023 56355
rect 36737 56321 36771 56355
rect 37289 56321 37323 56355
rect 39129 56321 39163 56355
rect 39589 56321 39623 56355
rect 40233 56321 40267 56355
rect 41521 56321 41555 56355
rect 43637 56321 43671 56355
rect 45293 56321 45327 56355
rect 49985 56321 50019 56355
rect 50813 56321 50847 56355
rect 52101 56321 52135 56355
rect 52377 56321 52411 56355
rect 53113 56321 53147 56355
rect 53573 56321 53607 56355
rect 54217 56321 54251 56355
rect 15117 56253 15151 56287
rect 16313 56253 16347 56287
rect 18061 56253 18095 56287
rect 18705 56253 18739 56287
rect 18797 56253 18831 56287
rect 19257 56253 19291 56287
rect 19349 56253 19383 56287
rect 21649 56253 21683 56287
rect 22017 56253 22051 56287
rect 22109 56253 22143 56287
rect 23305 56253 23339 56287
rect 24961 56253 24995 56287
rect 26157 56253 26191 56287
rect 27537 56253 27571 56287
rect 28733 56253 28767 56287
rect 28825 56253 28859 56287
rect 32689 56253 32723 56287
rect 34069 56253 34103 56287
rect 34253 56253 34287 56287
rect 36461 56253 36495 56287
rect 38209 56253 38243 56287
rect 40417 56253 40451 56287
rect 42901 56253 42935 56287
rect 42993 56253 43027 56287
rect 43729 56253 43763 56287
rect 43821 56253 43855 56287
rect 44189 56253 44223 56287
rect 44373 56253 44407 56287
rect 45477 56253 45511 56287
rect 49065 56253 49099 56287
rect 51181 56253 51215 56287
rect 53297 56253 53331 56287
rect 17233 56185 17267 56219
rect 22569 56185 22603 56219
rect 25605 56185 25639 56219
rect 37105 56185 37139 56219
rect 38853 56185 38887 56219
rect 39865 56185 39899 56219
rect 49709 56185 49743 56219
rect 50997 56185 51031 56219
rect 51825 56185 51859 56219
rect 15669 56117 15703 56151
rect 15761 56117 15795 56151
rect 17417 56117 17451 56151
rect 18245 56117 18279 56151
rect 19809 56117 19843 56151
rect 19901 56117 19935 56151
rect 22661 56117 22695 56151
rect 24041 56117 24075 56151
rect 25697 56117 25731 56151
rect 26985 56117 27019 56151
rect 28273 56117 28307 56151
rect 31953 56117 31987 56151
rect 34805 56117 34839 56151
rect 37473 56117 37507 56151
rect 38945 56117 38979 56151
rect 39773 56117 39807 56151
rect 41705 56117 41739 56151
rect 43269 56117 43303 56151
rect 44833 56117 44867 56151
rect 44925 56117 44959 56151
rect 51917 56117 51951 56151
rect 52193 56117 52227 56151
rect 16589 55913 16623 55947
rect 18153 55913 18187 55947
rect 20900 55913 20934 55947
rect 43637 55913 43671 55947
rect 45017 55913 45051 55947
rect 53113 55913 53147 55947
rect 16221 55845 16255 55879
rect 18521 55845 18555 55879
rect 24225 55845 24259 55879
rect 27997 55845 28031 55879
rect 29561 55845 29595 55879
rect 17141 55777 17175 55811
rect 17601 55777 17635 55811
rect 17693 55777 17727 55811
rect 20637 55777 20671 55811
rect 22477 55777 22511 55811
rect 26525 55777 26559 55811
rect 30113 55777 30147 55811
rect 51641 55777 51675 55811
rect 15761 55709 15795 55743
rect 16037 55709 16071 55743
rect 16313 55709 16347 55743
rect 17785 55709 17819 55743
rect 18337 55709 18371 55743
rect 18889 55709 18923 55743
rect 19257 55709 19291 55743
rect 19441 55709 19475 55743
rect 19717 55709 19751 55743
rect 26249 55709 26283 55743
rect 28089 55709 28123 55743
rect 35541 55709 35575 55743
rect 43453 55709 43487 55743
rect 44189 55709 44223 55743
rect 44373 55709 44407 55743
rect 44833 55709 44867 55743
rect 45569 55709 45603 55743
rect 51365 55709 51399 55743
rect 19625 55641 19659 55675
rect 22753 55641 22787 55675
rect 24777 55641 24811 55675
rect 36277 55641 36311 55675
rect 38025 55641 38059 55675
rect 15945 55573 15979 55607
rect 16497 55573 16531 55607
rect 16957 55573 16991 55607
rect 17049 55573 17083 55607
rect 19073 55573 19107 55607
rect 19901 55573 19935 55607
rect 22385 55573 22419 55607
rect 24501 55573 24535 55607
rect 28273 55573 28307 55607
rect 35449 55573 35483 55607
rect 43269 55573 43303 55607
rect 44557 55573 44591 55607
rect 44649 55573 44683 55607
rect 17693 55369 17727 55403
rect 19901 55369 19935 55403
rect 26525 55369 26559 55403
rect 29929 55369 29963 55403
rect 35725 55369 35759 55403
rect 39773 55369 39807 55403
rect 41613 55369 41647 55403
rect 44741 55369 44775 55403
rect 54493 55369 54527 55403
rect 25053 55301 25087 55335
rect 28457 55301 28491 55335
rect 32413 55301 32447 55335
rect 43269 55301 43303 55335
rect 51089 55301 51123 55335
rect 17141 55233 17175 55267
rect 17509 55233 17543 55267
rect 19809 55233 19843 55267
rect 21649 55233 21683 55267
rect 22477 55233 22511 55267
rect 24685 55233 24719 55267
rect 28181 55233 28215 55267
rect 32137 55233 32171 55267
rect 33977 55233 34011 55267
rect 39865 55233 39899 55267
rect 44833 55233 44867 55267
rect 48881 55233 48915 55267
rect 50813 55233 50847 55267
rect 52745 55233 52779 55267
rect 16957 55165 16991 55199
rect 18061 55165 18095 55199
rect 19533 55165 19567 55199
rect 21373 55165 21407 55199
rect 21833 55165 21867 55199
rect 22937 55165 22971 55199
rect 24409 55165 24443 55199
rect 24777 55165 24811 55199
rect 34253 55165 34287 55199
rect 38025 55165 38059 55199
rect 40141 55165 40175 55199
rect 42993 55165 43027 55199
rect 45109 55165 45143 55199
rect 46581 55165 46615 55199
rect 49157 55165 49191 55199
rect 50629 55165 50663 55199
rect 52561 55165 52595 55199
rect 53021 55165 53055 55199
rect 33885 55029 33919 55063
rect 38288 55029 38322 55063
rect 20637 54825 20671 54859
rect 24225 54825 24259 54859
rect 29377 54825 29411 54859
rect 36277 54825 36311 54859
rect 41153 54825 41187 54859
rect 43453 54825 43487 54859
rect 53113 54825 53147 54859
rect 26249 54757 26283 54791
rect 22385 54689 22419 54723
rect 22477 54689 22511 54723
rect 22753 54689 22787 54723
rect 27629 54689 27663 54723
rect 27905 54689 27939 54723
rect 37749 54689 37783 54723
rect 38025 54689 38059 54723
rect 41705 54689 41739 54723
rect 46765 54689 46799 54723
rect 51365 54689 51399 54723
rect 51641 54689 51675 54723
rect 53573 54621 53607 54655
rect 22109 54553 22143 54587
rect 27537 54553 27571 54587
rect 39865 54553 39899 54587
rect 41981 54553 42015 54587
rect 45017 54553 45051 54587
rect 53205 54553 53239 54587
rect 44373 54213 44407 54247
rect 44097 54145 44131 54179
rect 21373 54077 21407 54111
rect 21649 54077 21683 54111
rect 45845 54077 45879 54111
rect 19901 53941 19935 53975
rect 20729 53737 20763 53771
rect 26525 53737 26559 53771
rect 22477 53601 22511 53635
rect 27813 53533 27847 53567
rect 22201 53465 22235 53499
rect 19625 53193 19659 53227
rect 21373 53057 21407 53091
rect 21097 52989 21131 53023
rect 58265 44897 58299 44931
rect 58541 44829 58575 44863
<< metal1 >>
rect 1104 57690 58880 57712
rect 1104 57638 3010 57690
rect 3062 57638 3074 57690
rect 3126 57638 3138 57690
rect 3190 57638 3202 57690
rect 3254 57638 3266 57690
rect 3318 57638 33730 57690
rect 33782 57638 33794 57690
rect 33846 57638 33858 57690
rect 33910 57638 33922 57690
rect 33974 57638 33986 57690
rect 34038 57638 58880 57690
rect 1104 57616 58880 57638
rect 6730 57536 6736 57588
rect 6788 57576 6794 57588
rect 6917 57579 6975 57585
rect 6917 57576 6929 57579
rect 6788 57548 6929 57576
rect 6788 57536 6794 57548
rect 6917 57545 6929 57548
rect 6963 57545 6975 57579
rect 15286 57576 15292 57588
rect 6917 57539 6975 57545
rect 11072 57548 15292 57576
rect 2866 57468 2872 57520
rect 2924 57508 2930 57520
rect 2961 57511 3019 57517
rect 2961 57508 2973 57511
rect 2924 57480 2973 57508
rect 2924 57468 2930 57480
rect 2961 57477 2973 57480
rect 3007 57477 3019 57511
rect 2961 57471 3019 57477
rect 4798 57468 4804 57520
rect 4856 57508 4862 57520
rect 4893 57511 4951 57517
rect 4893 57508 4905 57511
rect 4856 57480 4905 57508
rect 4856 57468 4862 57480
rect 4893 57477 4905 57480
rect 4939 57477 4951 57511
rect 4893 57471 4951 57477
rect 8662 57468 8668 57520
rect 8720 57508 8726 57520
rect 8941 57511 8999 57517
rect 8941 57508 8953 57511
rect 8720 57480 8953 57508
rect 8720 57468 8726 57480
rect 8941 57477 8953 57480
rect 8987 57477 8999 57511
rect 8941 57471 8999 57477
rect 10594 57468 10600 57520
rect 10652 57508 10658 57520
rect 11072 57517 11100 57548
rect 15286 57536 15292 57548
rect 15344 57536 15350 57588
rect 26234 57536 26240 57588
rect 26292 57536 26298 57588
rect 27982 57536 27988 57588
rect 28040 57576 28046 57588
rect 28261 57579 28319 57585
rect 28261 57576 28273 57579
rect 28040 57548 28273 57576
rect 28040 57536 28046 57548
rect 28261 57545 28273 57548
rect 28307 57545 28319 57579
rect 28261 57539 28319 57545
rect 30374 57536 30380 57588
rect 30432 57536 30438 57588
rect 34146 57536 34152 57588
rect 34204 57536 34210 57588
rect 35710 57536 35716 57588
rect 35768 57576 35774 57588
rect 35897 57579 35955 57585
rect 35897 57576 35909 57579
rect 35768 57548 35909 57576
rect 35768 57536 35774 57548
rect 35897 57545 35909 57548
rect 35943 57545 35955 57579
rect 35897 57539 35955 57545
rect 45370 57536 45376 57588
rect 45428 57576 45434 57588
rect 45649 57579 45707 57585
rect 45649 57576 45661 57579
rect 45428 57548 45661 57576
rect 45428 57536 45434 57548
rect 45649 57545 45661 57548
rect 45695 57545 45707 57579
rect 45649 57539 45707 57545
rect 47302 57536 47308 57588
rect 47360 57576 47366 57588
rect 47765 57579 47823 57585
rect 47765 57576 47777 57579
rect 47360 57548 47777 57576
rect 47360 57536 47366 57548
rect 47765 57545 47777 57548
rect 47811 57545 47823 57579
rect 47765 57539 47823 57545
rect 49694 57536 49700 57588
rect 49752 57536 49758 57588
rect 51166 57536 51172 57588
rect 51224 57576 51230 57588
rect 51445 57579 51503 57585
rect 51445 57576 51457 57579
rect 51224 57548 51457 57576
rect 51224 57536 51230 57548
rect 51445 57545 51457 57548
rect 51491 57545 51503 57579
rect 51445 57539 51503 57545
rect 53098 57536 53104 57588
rect 53156 57576 53162 57588
rect 53377 57579 53435 57585
rect 53377 57576 53389 57579
rect 53156 57548 53389 57576
rect 53156 57536 53162 57548
rect 53377 57545 53389 57548
rect 53423 57545 53435 57579
rect 53377 57539 53435 57545
rect 55030 57536 55036 57588
rect 55088 57576 55094 57588
rect 55493 57579 55551 57585
rect 55493 57576 55505 57579
rect 55088 57548 55505 57576
rect 55088 57536 55094 57548
rect 55493 57545 55505 57548
rect 55539 57545 55551 57579
rect 55493 57539 55551 57545
rect 56962 57536 56968 57588
rect 57020 57576 57026 57588
rect 57241 57579 57299 57585
rect 57241 57576 57253 57579
rect 57020 57548 57253 57576
rect 57020 57536 57026 57548
rect 57241 57545 57253 57548
rect 57287 57545 57299 57579
rect 57241 57539 57299 57545
rect 10689 57511 10747 57517
rect 10689 57508 10701 57511
rect 10652 57480 10701 57508
rect 10652 57468 10658 57480
rect 10689 57477 10701 57480
rect 10735 57477 10747 57511
rect 10689 57471 10747 57477
rect 11057 57511 11115 57517
rect 11057 57477 11069 57511
rect 11103 57477 11115 57511
rect 11057 57471 11115 57477
rect 12526 57468 12532 57520
rect 12584 57508 12590 57520
rect 12621 57511 12679 57517
rect 12621 57508 12633 57511
rect 12584 57480 12633 57508
rect 12584 57468 12590 57480
rect 12621 57477 12633 57480
rect 12667 57477 12679 57511
rect 12621 57471 12679 57477
rect 12912 57480 14412 57508
rect 934 57400 940 57452
rect 992 57440 998 57452
rect 1397 57443 1455 57449
rect 1397 57440 1409 57443
rect 992 57412 1409 57440
rect 992 57400 998 57412
rect 1397 57409 1409 57412
rect 1443 57409 1455 57443
rect 1397 57403 1455 57409
rect 3329 57443 3387 57449
rect 3329 57409 3341 57443
rect 3375 57440 3387 57443
rect 4062 57440 4068 57452
rect 3375 57412 4068 57440
rect 3375 57409 3387 57412
rect 3329 57403 3387 57409
rect 4062 57400 4068 57412
rect 4120 57400 4126 57452
rect 5258 57400 5264 57452
rect 5316 57400 5322 57452
rect 7190 57400 7196 57452
rect 7248 57400 7254 57452
rect 9309 57443 9367 57449
rect 9309 57409 9321 57443
rect 9355 57440 9367 57443
rect 12912 57440 12940 57480
rect 9355 57412 12940 57440
rect 12989 57443 13047 57449
rect 9355 57409 9367 57412
rect 9309 57403 9367 57409
rect 12989 57409 13001 57443
rect 13035 57409 13047 57443
rect 14384 57440 14412 57480
rect 14458 57468 14464 57520
rect 14516 57508 14522 57520
rect 14553 57511 14611 57517
rect 14553 57508 14565 57511
rect 14516 57480 14565 57508
rect 14516 57468 14522 57480
rect 14553 57477 14565 57480
rect 14599 57477 14611 57511
rect 15194 57508 15200 57520
rect 14553 57471 14611 57477
rect 14844 57480 15200 57508
rect 14844 57440 14872 57480
rect 15194 57468 15200 57480
rect 15252 57468 15258 57520
rect 16390 57468 16396 57520
rect 16448 57508 16454 57520
rect 16669 57511 16727 57517
rect 16669 57508 16681 57511
rect 16448 57480 16681 57508
rect 16448 57468 16454 57480
rect 16669 57477 16681 57480
rect 16715 57477 16727 57511
rect 16669 57471 16727 57477
rect 18322 57468 18328 57520
rect 18380 57508 18386 57520
rect 18417 57511 18475 57517
rect 18417 57508 18429 57511
rect 18380 57480 18429 57508
rect 18380 57468 18386 57480
rect 18417 57477 18429 57480
rect 18463 57477 18475 57511
rect 18417 57471 18475 57477
rect 20254 57468 20260 57520
rect 20312 57508 20318 57520
rect 20349 57511 20407 57517
rect 20349 57508 20361 57511
rect 20312 57480 20361 57508
rect 20312 57468 20318 57480
rect 20349 57477 20361 57480
rect 20395 57477 20407 57511
rect 20349 57471 20407 57477
rect 22186 57468 22192 57520
rect 22244 57508 22250 57520
rect 22281 57511 22339 57517
rect 22281 57508 22293 57511
rect 22244 57480 22293 57508
rect 22244 57468 22250 57480
rect 22281 57477 22293 57480
rect 22327 57477 22339 57511
rect 22281 57471 22339 57477
rect 24118 57468 24124 57520
rect 24176 57508 24182 57520
rect 24397 57511 24455 57517
rect 24397 57508 24409 57511
rect 24176 57480 24409 57508
rect 24176 57468 24182 57480
rect 24397 57477 24409 57480
rect 24443 57477 24455 57511
rect 24397 57471 24455 57477
rect 31846 57468 31852 57520
rect 31904 57508 31910 57520
rect 32125 57511 32183 57517
rect 32125 57508 32137 57511
rect 31904 57480 32137 57508
rect 31904 57468 31910 57480
rect 32125 57477 32137 57480
rect 32171 57477 32183 57511
rect 32125 57471 32183 57477
rect 37642 57468 37648 57520
rect 37700 57508 37706 57520
rect 37737 57511 37795 57517
rect 37737 57508 37749 57511
rect 37700 57480 37749 57508
rect 37700 57468 37706 57480
rect 37737 57477 37749 57480
rect 37783 57477 37795 57511
rect 37737 57471 37795 57477
rect 39574 57468 39580 57520
rect 39632 57508 39638 57520
rect 39853 57511 39911 57517
rect 39853 57508 39865 57511
rect 39632 57480 39865 57508
rect 39632 57468 39638 57480
rect 39853 57477 39865 57480
rect 39899 57477 39911 57511
rect 39853 57471 39911 57477
rect 41506 57468 41512 57520
rect 41564 57508 41570 57520
rect 41601 57511 41659 57517
rect 41601 57508 41613 57511
rect 41564 57480 41613 57508
rect 41564 57468 41570 57480
rect 41601 57477 41613 57480
rect 41647 57477 41659 57511
rect 41601 57471 41659 57477
rect 43438 57468 43444 57520
rect 43496 57508 43502 57520
rect 43533 57511 43591 57517
rect 43533 57508 43545 57511
rect 43496 57480 43545 57508
rect 43496 57468 43502 57480
rect 43533 57477 43545 57480
rect 43579 57477 43591 57511
rect 43533 57471 43591 57477
rect 53006 57468 53012 57520
rect 53064 57508 53070 57520
rect 55401 57511 55459 57517
rect 55401 57508 55413 57511
rect 53064 57480 55413 57508
rect 53064 57468 53070 57480
rect 55401 57477 55413 57480
rect 55447 57477 55459 57511
rect 55401 57471 55459 57477
rect 56134 57468 56140 57520
rect 56192 57508 56198 57520
rect 58161 57511 58219 57517
rect 58161 57508 58173 57511
rect 56192 57480 58173 57508
rect 56192 57468 56198 57480
rect 58161 57477 58173 57480
rect 58207 57477 58219 57511
rect 58161 57471 58219 57477
rect 58529 57511 58587 57517
rect 58529 57477 58541 57511
rect 58575 57508 58587 57511
rect 58894 57508 58900 57520
rect 58575 57480 58900 57508
rect 58575 57477 58587 57480
rect 58529 57471 58587 57477
rect 58894 57468 58900 57480
rect 58952 57468 58958 57520
rect 14384 57412 14872 57440
rect 14921 57443 14979 57449
rect 12989 57403 13047 57409
rect 14921 57409 14933 57443
rect 14967 57440 14979 57443
rect 16758 57440 16764 57452
rect 14967 57412 16764 57440
rect 14967 57409 14979 57412
rect 14921 57403 14979 57409
rect 1673 57375 1731 57381
rect 1673 57341 1685 57375
rect 1719 57372 1731 57375
rect 1719 57344 6914 57372
rect 1719 57341 1731 57344
rect 1673 57335 1731 57341
rect 6886 57236 6914 57344
rect 13004 57304 13032 57403
rect 16758 57400 16764 57412
rect 16816 57400 16822 57452
rect 17037 57443 17095 57449
rect 17037 57409 17049 57443
rect 17083 57440 17095 57443
rect 17218 57440 17224 57452
rect 17083 57412 17224 57440
rect 17083 57409 17095 57412
rect 17037 57403 17095 57409
rect 17218 57400 17224 57412
rect 17276 57400 17282 57452
rect 18785 57443 18843 57449
rect 18785 57409 18797 57443
rect 18831 57440 18843 57443
rect 18874 57440 18880 57452
rect 18831 57412 18880 57440
rect 18831 57409 18843 57412
rect 18785 57403 18843 57409
rect 18874 57400 18880 57412
rect 18932 57400 18938 57452
rect 20714 57400 20720 57452
rect 20772 57400 20778 57452
rect 22462 57400 22468 57452
rect 22520 57440 22526 57452
rect 22649 57443 22707 57449
rect 22649 57440 22661 57443
rect 22520 57412 22661 57440
rect 22520 57400 22526 57412
rect 22649 57409 22661 57412
rect 22695 57409 22707 57443
rect 22649 57403 22707 57409
rect 24762 57400 24768 57452
rect 24820 57400 24826 57452
rect 26513 57443 26571 57449
rect 26513 57409 26525 57443
rect 26559 57440 26571 57443
rect 27062 57440 27068 57452
rect 26559 57412 27068 57440
rect 26559 57409 26571 57412
rect 26513 57403 26571 57409
rect 27062 57400 27068 57412
rect 27120 57400 27126 57452
rect 27706 57400 27712 57452
rect 27764 57440 27770 57452
rect 28169 57443 28227 57449
rect 28169 57440 28181 57443
rect 27764 57412 28181 57440
rect 27764 57400 27770 57412
rect 28169 57409 28181 57412
rect 28215 57409 28227 57443
rect 28169 57403 28227 57409
rect 30098 57400 30104 57452
rect 30156 57400 30162 57452
rect 32490 57400 32496 57452
rect 32548 57400 32554 57452
rect 34238 57400 34244 57452
rect 34296 57400 34302 57452
rect 35894 57400 35900 57452
rect 35952 57440 35958 57452
rect 36173 57443 36231 57449
rect 36173 57440 36185 57443
rect 35952 57412 36185 57440
rect 35952 57400 35958 57412
rect 36173 57409 36185 57412
rect 36219 57409 36231 57443
rect 36173 57403 36231 57409
rect 38102 57400 38108 57452
rect 38160 57400 38166 57452
rect 40218 57400 40224 57452
rect 40276 57400 40282 57452
rect 41966 57400 41972 57452
rect 42024 57400 42030 57452
rect 43898 57400 43904 57452
rect 43956 57400 43962 57452
rect 45554 57400 45560 57452
rect 45612 57400 45618 57452
rect 47670 57400 47676 57452
rect 47728 57400 47734 57452
rect 49418 57400 49424 57452
rect 49476 57400 49482 57452
rect 51166 57400 51172 57452
rect 51224 57440 51230 57452
rect 51353 57443 51411 57449
rect 51353 57440 51365 57443
rect 51224 57412 51365 57440
rect 51224 57400 51230 57412
rect 51353 57409 51365 57412
rect 51399 57409 51411 57443
rect 51353 57403 51411 57409
rect 51994 57400 52000 57452
rect 52052 57440 52058 57452
rect 53285 57443 53343 57449
rect 53285 57440 53297 57443
rect 52052 57412 53297 57440
rect 52052 57400 52058 57412
rect 53285 57409 53297 57412
rect 53331 57409 53343 57443
rect 53285 57403 53343 57409
rect 55858 57400 55864 57452
rect 55916 57440 55922 57452
rect 57149 57443 57207 57449
rect 57149 57440 57161 57443
rect 55916 57412 57161 57440
rect 55916 57400 55922 57412
rect 57149 57409 57161 57412
rect 57195 57409 57207 57443
rect 57149 57403 57207 57409
rect 16850 57372 16856 57384
rect 16546 57344 16856 57372
rect 16114 57304 16120 57316
rect 13004 57276 16120 57304
rect 16114 57264 16120 57276
rect 16172 57264 16178 57316
rect 16546 57236 16574 57344
rect 16850 57332 16856 57344
rect 16908 57332 16914 57384
rect 6886 57208 16574 57236
rect 1104 57146 58880 57168
rect 1104 57094 2350 57146
rect 2402 57094 2414 57146
rect 2466 57094 2478 57146
rect 2530 57094 2542 57146
rect 2594 57094 2606 57146
rect 2658 57094 33070 57146
rect 33122 57094 33134 57146
rect 33186 57094 33198 57146
rect 33250 57094 33262 57146
rect 33314 57094 33326 57146
rect 33378 57094 58880 57146
rect 1104 57072 58880 57094
rect 6886 57004 15976 57032
rect 5258 56924 5264 56976
rect 5316 56964 5322 56976
rect 6886 56964 6914 57004
rect 5316 56936 6914 56964
rect 15841 56967 15899 56973
rect 5316 56924 5322 56936
rect 15841 56933 15853 56967
rect 15887 56933 15899 56967
rect 15948 56964 15976 57004
rect 16022 56992 16028 57044
rect 16080 57032 16086 57044
rect 16853 57035 16911 57041
rect 16080 57004 16804 57032
rect 16080 56992 16086 57004
rect 16776 56964 16804 57004
rect 16853 57001 16865 57035
rect 16899 57032 16911 57035
rect 21266 57032 21272 57044
rect 16899 57004 21272 57032
rect 16899 57001 16911 57004
rect 16853 56995 16911 57001
rect 21266 56992 21272 57004
rect 21324 56992 21330 57044
rect 51534 56992 51540 57044
rect 51592 57032 51598 57044
rect 52270 57032 52276 57044
rect 51592 57004 52276 57032
rect 51592 56992 51598 57004
rect 52270 56992 52276 57004
rect 52328 57032 52334 57044
rect 52328 57004 52960 57032
rect 52328 56992 52334 57004
rect 20806 56964 20812 56976
rect 15948 56936 16574 56964
rect 16776 56936 20812 56964
rect 15841 56927 15899 56933
rect 15565 56831 15623 56837
rect 15565 56797 15577 56831
rect 15611 56828 15623 56831
rect 15856 56828 15884 56927
rect 16390 56856 16396 56908
rect 16448 56856 16454 56908
rect 16546 56896 16574 56936
rect 20806 56924 20812 56936
rect 20864 56924 20870 56976
rect 51074 56924 51080 56976
rect 51132 56964 51138 56976
rect 52549 56967 52607 56973
rect 52549 56964 52561 56967
rect 51132 56936 52561 56964
rect 51132 56924 51138 56936
rect 52549 56933 52561 56936
rect 52595 56933 52607 56967
rect 52932 56964 52960 57004
rect 52932 56936 53144 56964
rect 52549 56927 52607 56933
rect 17126 56896 17132 56908
rect 16546 56868 17132 56896
rect 17126 56856 17132 56868
rect 17184 56856 17190 56908
rect 17310 56856 17316 56908
rect 17368 56896 17374 56908
rect 17497 56899 17555 56905
rect 17497 56896 17509 56899
rect 17368 56868 17509 56896
rect 17368 56856 17374 56868
rect 17497 56865 17509 56868
rect 17543 56865 17555 56899
rect 17497 56859 17555 56865
rect 17862 56856 17868 56908
rect 17920 56896 17926 56908
rect 21913 56899 21971 56905
rect 21913 56896 21925 56899
rect 17920 56868 21925 56896
rect 17920 56856 17926 56868
rect 21913 56865 21925 56868
rect 21959 56865 21971 56899
rect 21913 56859 21971 56865
rect 51534 56856 51540 56908
rect 51592 56896 51598 56908
rect 51813 56899 51871 56905
rect 51813 56896 51825 56899
rect 51592 56868 51825 56896
rect 51592 56856 51598 56868
rect 51813 56865 51825 56868
rect 51859 56865 51871 56899
rect 51813 56859 51871 56865
rect 51994 56856 52000 56908
rect 52052 56856 52058 56908
rect 53006 56856 53012 56908
rect 53064 56856 53070 56908
rect 53116 56905 53144 56936
rect 53101 56899 53159 56905
rect 53101 56865 53113 56899
rect 53147 56865 53159 56899
rect 53101 56859 53159 56865
rect 15611 56800 15884 56828
rect 15611 56797 15623 56800
rect 15565 56791 15623 56797
rect 15930 56788 15936 56840
rect 15988 56828 15994 56840
rect 16206 56828 16212 56840
rect 15988 56800 16212 56828
rect 15988 56788 15994 56800
rect 16206 56788 16212 56800
rect 16264 56788 16270 56840
rect 16666 56788 16672 56840
rect 16724 56788 16730 56840
rect 16850 56788 16856 56840
rect 16908 56828 16914 56840
rect 17773 56831 17831 56837
rect 17773 56828 17785 56831
rect 16908 56800 17785 56828
rect 16908 56788 16914 56800
rect 17773 56797 17785 56800
rect 17819 56797 17831 56831
rect 17773 56791 17831 56797
rect 18138 56788 18144 56840
rect 18196 56828 18202 56840
rect 18325 56831 18383 56837
rect 18325 56828 18337 56831
rect 18196 56800 18337 56828
rect 18196 56788 18202 56800
rect 18325 56797 18337 56800
rect 18371 56797 18383 56831
rect 19518 56828 19524 56840
rect 18325 56791 18383 56797
rect 18432 56800 19524 56828
rect 7190 56720 7196 56772
rect 7248 56760 7254 56772
rect 16301 56763 16359 56769
rect 16301 56760 16313 56763
rect 7248 56732 16313 56760
rect 7248 56720 7254 56732
rect 16301 56729 16313 56732
rect 16347 56760 16359 56763
rect 17313 56763 17371 56769
rect 17313 56760 17325 56763
rect 16347 56732 17325 56760
rect 16347 56729 16359 56732
rect 16301 56723 16359 56729
rect 17313 56729 17325 56732
rect 17359 56760 17371 56763
rect 17954 56760 17960 56772
rect 17359 56732 17960 56760
rect 17359 56729 17371 56732
rect 17313 56723 17371 56729
rect 17954 56720 17960 56732
rect 18012 56720 18018 56772
rect 18049 56763 18107 56769
rect 18049 56729 18061 56763
rect 18095 56760 18107 56763
rect 18432 56760 18460 56800
rect 19518 56788 19524 56800
rect 19576 56788 19582 56840
rect 22186 56788 22192 56840
rect 22244 56788 22250 56840
rect 22462 56788 22468 56840
rect 22520 56828 22526 56840
rect 23017 56831 23075 56837
rect 23017 56828 23029 56831
rect 22520 56800 23029 56828
rect 22520 56788 22526 56800
rect 23017 56797 23029 56800
rect 23063 56797 23075 56831
rect 23017 56791 23075 56797
rect 27062 56788 27068 56840
rect 27120 56788 27126 56840
rect 27798 56788 27804 56840
rect 27856 56788 27862 56840
rect 28166 56788 28172 56840
rect 28224 56788 28230 56840
rect 51445 56831 51503 56837
rect 51445 56797 51457 56831
rect 51491 56828 51503 56831
rect 52730 56828 52736 56840
rect 51491 56800 52736 56828
rect 51491 56797 51503 56800
rect 51445 56791 51503 56797
rect 52730 56788 52736 56800
rect 52788 56788 52794 56840
rect 18095 56732 18460 56760
rect 18524 56732 20668 56760
rect 18095 56729 18107 56732
rect 18049 56723 18107 56729
rect 15749 56695 15807 56701
rect 15749 56661 15761 56695
rect 15795 56692 15807 56695
rect 16022 56692 16028 56704
rect 15795 56664 16028 56692
rect 15795 56661 15807 56664
rect 15749 56655 15807 56661
rect 16022 56652 16028 56664
rect 16080 56652 16086 56704
rect 16942 56652 16948 56704
rect 17000 56652 17006 56704
rect 17126 56652 17132 56704
rect 17184 56692 17190 56704
rect 17402 56692 17408 56704
rect 17184 56664 17408 56692
rect 17184 56652 17190 56664
rect 17402 56652 17408 56664
rect 17460 56652 17466 56704
rect 18524 56701 18552 56732
rect 18509 56695 18567 56701
rect 18509 56661 18521 56695
rect 18555 56661 18567 56695
rect 18509 56655 18567 56661
rect 18598 56652 18604 56704
rect 18656 56692 18662 56704
rect 20441 56695 20499 56701
rect 20441 56692 20453 56695
rect 18656 56664 20453 56692
rect 18656 56652 18662 56664
rect 20441 56661 20453 56664
rect 20487 56661 20499 56695
rect 20640 56692 20668 56732
rect 20898 56720 20904 56772
rect 20956 56720 20962 56772
rect 52089 56763 52147 56769
rect 52089 56729 52101 56763
rect 52135 56760 52147 56763
rect 53024 56760 53052 56856
rect 52135 56732 53052 56760
rect 52135 56729 52147 56732
rect 52089 56723 52147 56729
rect 22554 56692 22560 56704
rect 20640 56664 22560 56692
rect 20441 56655 20499 56661
rect 22554 56652 22560 56664
rect 22612 56652 22618 56704
rect 23658 56652 23664 56704
rect 23716 56652 23722 56704
rect 26510 56652 26516 56704
rect 26568 56652 26574 56704
rect 27154 56652 27160 56704
rect 27212 56692 27218 56704
rect 27249 56695 27307 56701
rect 27249 56692 27261 56695
rect 27212 56664 27261 56692
rect 27212 56652 27218 56664
rect 27249 56661 27261 56664
rect 27295 56661 27307 56695
rect 27249 56655 27307 56661
rect 27890 56652 27896 56704
rect 27948 56692 27954 56704
rect 27985 56695 28043 56701
rect 27985 56692 27997 56695
rect 27948 56664 27997 56692
rect 27948 56652 27954 56664
rect 27985 56661 27997 56664
rect 28031 56661 28043 56695
rect 27985 56655 28043 56661
rect 51626 56652 51632 56704
rect 51684 56652 51690 56704
rect 52454 56652 52460 56704
rect 52512 56652 52518 56704
rect 52914 56652 52920 56704
rect 52972 56652 52978 56704
rect 1104 56602 58880 56624
rect 1104 56550 3010 56602
rect 3062 56550 3074 56602
rect 3126 56550 3138 56602
rect 3190 56550 3202 56602
rect 3254 56550 3266 56602
rect 3318 56550 33730 56602
rect 33782 56550 33794 56602
rect 33846 56550 33858 56602
rect 33910 56550 33922 56602
rect 33974 56550 33986 56602
rect 34038 56550 58880 56602
rect 1104 56528 58880 56550
rect 15194 56448 15200 56500
rect 15252 56448 15258 56500
rect 15286 56448 15292 56500
rect 15344 56488 15350 56500
rect 16209 56491 16267 56497
rect 16209 56488 16221 56491
rect 15344 56460 16221 56488
rect 15344 56448 15350 56460
rect 16209 56457 16221 56460
rect 16255 56488 16267 56491
rect 16255 56460 16712 56488
rect 16255 56457 16267 56460
rect 16209 56451 16267 56457
rect 15212 56420 15240 56448
rect 15930 56420 15936 56432
rect 15212 56392 15936 56420
rect 15930 56380 15936 56392
rect 15988 56380 15994 56432
rect 16114 56380 16120 56432
rect 16172 56380 16178 56432
rect 16684 56352 16712 56460
rect 16758 56448 16764 56500
rect 16816 56488 16822 56500
rect 17770 56488 17776 56500
rect 16816 56460 17776 56488
rect 16816 56448 16822 56460
rect 17770 56448 17776 56460
rect 17828 56488 17834 56500
rect 17865 56491 17923 56497
rect 17865 56488 17877 56491
rect 17828 56460 17877 56488
rect 17828 56448 17834 56460
rect 17865 56457 17877 56460
rect 17911 56457 17923 56491
rect 19242 56488 19248 56500
rect 17865 56451 17923 56457
rect 17972 56460 19248 56488
rect 16850 56380 16856 56432
rect 16908 56420 16914 56432
rect 16945 56423 17003 56429
rect 16945 56420 16957 56423
rect 16908 56392 16957 56420
rect 16908 56380 16914 56392
rect 16945 56389 16957 56392
rect 16991 56389 17003 56423
rect 17972 56420 18000 56460
rect 19242 56448 19248 56460
rect 19300 56448 19306 56500
rect 23477 56491 23535 56497
rect 19352 56460 22048 56488
rect 19352 56420 19380 56460
rect 16945 56383 17003 56389
rect 17144 56392 18000 56420
rect 19260 56392 19380 56420
rect 17144 56356 17172 56392
rect 17052 56352 17172 56356
rect 16684 56328 17172 56352
rect 16684 56324 17080 56328
rect 17218 56312 17224 56364
rect 17276 56352 17282 56364
rect 17773 56355 17831 56361
rect 17773 56352 17785 56355
rect 17276 56324 17785 56352
rect 17276 56312 17282 56324
rect 17773 56321 17785 56324
rect 17819 56352 17831 56355
rect 18601 56355 18659 56361
rect 17819 56324 18276 56352
rect 17819 56321 17831 56324
rect 17773 56315 17831 56321
rect 15105 56287 15163 56293
rect 15105 56253 15117 56287
rect 15151 56253 15163 56287
rect 15105 56247 15163 56253
rect 16301 56287 16359 56293
rect 16301 56253 16313 56287
rect 16347 56284 16359 56287
rect 16390 56284 16396 56296
rect 16347 56256 16396 56284
rect 16347 56253 16359 56256
rect 16301 56247 16359 56253
rect 15120 56216 15148 56247
rect 16316 56216 16344 56247
rect 16390 56244 16396 56256
rect 16448 56284 16454 56296
rect 17310 56284 17316 56296
rect 16448 56256 17316 56284
rect 16448 56244 16454 56256
rect 17310 56244 17316 56256
rect 17368 56244 17374 56296
rect 18049 56287 18107 56293
rect 18049 56253 18061 56287
rect 18095 56253 18107 56287
rect 18248 56284 18276 56324
rect 18601 56321 18613 56355
rect 18647 56352 18659 56355
rect 18874 56352 18880 56364
rect 18647 56324 18880 56352
rect 18647 56321 18659 56324
rect 18601 56315 18659 56321
rect 18874 56312 18880 56324
rect 18932 56312 18938 56364
rect 18690 56284 18696 56296
rect 18248 56256 18696 56284
rect 18049 56247 18107 56253
rect 15120 56188 16344 56216
rect 17221 56219 17279 56225
rect 17221 56185 17233 56219
rect 17267 56216 17279 56219
rect 17586 56216 17592 56228
rect 17267 56188 17592 56216
rect 17267 56185 17279 56188
rect 17221 56179 17279 56185
rect 17586 56176 17592 56188
rect 17644 56216 17650 56228
rect 18064 56216 18092 56247
rect 18690 56244 18696 56256
rect 18748 56244 18754 56296
rect 19260 56293 19288 56392
rect 20898 56380 20904 56432
rect 20956 56380 20962 56432
rect 21266 56380 21272 56432
rect 21324 56420 21330 56432
rect 21361 56423 21419 56429
rect 21361 56420 21373 56423
rect 21324 56392 21373 56420
rect 21324 56380 21330 56392
rect 21361 56389 21373 56392
rect 21407 56389 21419 56423
rect 21361 56383 21419 56389
rect 22020 56420 22048 56460
rect 23477 56457 23489 56491
rect 23523 56488 23535 56491
rect 23658 56488 23664 56500
rect 23523 56460 23664 56488
rect 23523 56457 23535 56460
rect 23477 56451 23535 56457
rect 23658 56448 23664 56460
rect 23716 56448 23722 56500
rect 23937 56491 23995 56497
rect 23937 56457 23949 56491
rect 23983 56457 23995 56491
rect 23937 56451 23995 56457
rect 23569 56423 23627 56429
rect 22020 56392 23336 56420
rect 19426 56312 19432 56364
rect 19484 56312 19490 56364
rect 18785 56287 18843 56293
rect 18785 56253 18797 56287
rect 18831 56284 18843 56287
rect 19245 56287 19303 56293
rect 19245 56284 19257 56287
rect 18831 56256 19257 56284
rect 18831 56253 18843 56256
rect 18785 56247 18843 56253
rect 19245 56253 19257 56256
rect 19291 56253 19303 56287
rect 19245 56247 19303 56253
rect 19337 56287 19395 56293
rect 19337 56253 19349 56287
rect 19383 56284 19395 56287
rect 19978 56284 19984 56296
rect 19383 56256 19984 56284
rect 19383 56253 19395 56256
rect 19337 56247 19395 56253
rect 18800 56216 18828 56247
rect 17644 56188 18828 56216
rect 17644 56176 17650 56188
rect 18874 56176 18880 56228
rect 18932 56216 18938 56228
rect 19352 56216 19380 56247
rect 19978 56244 19984 56256
rect 20036 56244 20042 56296
rect 22020 56293 22048 56392
rect 22189 56355 22247 56361
rect 22189 56321 22201 56355
rect 22235 56352 22247 56355
rect 22462 56352 22468 56364
rect 22235 56324 22468 56352
rect 22235 56321 22247 56324
rect 22189 56315 22247 56321
rect 22462 56312 22468 56324
rect 22520 56312 22526 56364
rect 22833 56355 22891 56361
rect 22833 56352 22845 56355
rect 22572 56324 22845 56352
rect 21637 56287 21695 56293
rect 21637 56253 21649 56287
rect 21683 56253 21695 56287
rect 21637 56247 21695 56253
rect 22005 56287 22063 56293
rect 22005 56253 22017 56287
rect 22051 56253 22063 56287
rect 22005 56247 22063 56253
rect 22097 56287 22155 56293
rect 22097 56253 22109 56287
rect 22143 56284 22155 56287
rect 22278 56284 22284 56296
rect 22143 56256 22284 56284
rect 22143 56253 22155 56256
rect 22097 56247 22155 56253
rect 18932 56188 19380 56216
rect 18932 56176 18938 56188
rect 19426 56176 19432 56228
rect 19484 56216 19490 56228
rect 21652 56216 21680 56247
rect 22278 56244 22284 56256
rect 22336 56244 22342 56296
rect 22572 56225 22600 56324
rect 22833 56321 22845 56324
rect 22879 56321 22891 56355
rect 22833 56315 22891 56321
rect 23308 56293 23336 56392
rect 23569 56389 23581 56423
rect 23615 56420 23627 56423
rect 23750 56420 23756 56432
rect 23615 56392 23756 56420
rect 23615 56389 23627 56392
rect 23569 56383 23627 56389
rect 23750 56380 23756 56392
rect 23808 56380 23814 56432
rect 23952 56352 23980 56451
rect 24762 56448 24768 56500
rect 24820 56488 24826 56500
rect 25133 56491 25191 56497
rect 25133 56488 25145 56491
rect 24820 56460 25145 56488
rect 24820 56448 24826 56460
rect 25133 56457 25145 56460
rect 25179 56457 25191 56491
rect 26329 56491 26387 56497
rect 25133 56451 25191 56457
rect 25240 56460 26280 56488
rect 25240 56429 25268 56460
rect 25225 56423 25283 56429
rect 25225 56389 25237 56423
rect 25271 56389 25283 56423
rect 26252 56420 26280 56460
rect 26329 56457 26341 56491
rect 26375 56488 26387 56491
rect 26510 56488 26516 56500
rect 26375 56460 26516 56488
rect 26375 56457 26387 56460
rect 26329 56451 26387 56457
rect 26510 56448 26516 56460
rect 26568 56448 26574 56500
rect 26789 56491 26847 56497
rect 26789 56457 26801 56491
rect 26835 56488 26847 56491
rect 27798 56488 27804 56500
rect 26835 56460 27804 56488
rect 26835 56457 26847 56460
rect 26789 56451 26847 56457
rect 27798 56448 27804 56460
rect 27856 56448 27862 56500
rect 28166 56448 28172 56500
rect 28224 56448 28230 56500
rect 32125 56491 32183 56497
rect 32125 56457 32137 56491
rect 32171 56457 32183 56491
rect 32125 56451 32183 56457
rect 27062 56420 27068 56432
rect 25225 56383 25283 56389
rect 25792 56392 26188 56420
rect 26252 56392 27068 56420
rect 24213 56355 24271 56361
rect 24213 56352 24225 56355
rect 23952 56324 24225 56352
rect 24213 56321 24225 56324
rect 24259 56321 24271 56355
rect 25792 56352 25820 56392
rect 24213 56315 24271 56321
rect 24964 56324 25820 56352
rect 25869 56339 25927 56345
rect 24964 56293 24992 56324
rect 25869 56305 25881 56339
rect 25915 56305 25927 56339
rect 25869 56299 25927 56305
rect 23293 56287 23351 56293
rect 23293 56253 23305 56287
rect 23339 56253 23351 56287
rect 23293 56247 23351 56253
rect 24949 56287 25007 56293
rect 24949 56253 24961 56287
rect 24995 56253 25007 56287
rect 24949 56247 25007 56253
rect 22557 56219 22615 56225
rect 19484 56188 20024 56216
rect 21652 56188 22094 56216
rect 19484 56176 19490 56188
rect 15654 56108 15660 56160
rect 15712 56108 15718 56160
rect 15749 56151 15807 56157
rect 15749 56117 15761 56151
rect 15795 56148 15807 56151
rect 16022 56148 16028 56160
rect 15795 56120 16028 56148
rect 15795 56117 15807 56120
rect 15749 56111 15807 56117
rect 16022 56108 16028 56120
rect 16080 56108 16086 56160
rect 17405 56151 17463 56157
rect 17405 56117 17417 56151
rect 17451 56148 17463 56151
rect 17494 56148 17500 56160
rect 17451 56120 17500 56148
rect 17451 56117 17463 56120
rect 17405 56111 17463 56117
rect 17494 56108 17500 56120
rect 17552 56108 17558 56160
rect 18233 56151 18291 56157
rect 18233 56117 18245 56151
rect 18279 56148 18291 56151
rect 18322 56148 18328 56160
rect 18279 56120 18328 56148
rect 18279 56117 18291 56120
rect 18233 56111 18291 56117
rect 18322 56108 18328 56120
rect 18380 56108 18386 56160
rect 19334 56108 19340 56160
rect 19392 56148 19398 56160
rect 19610 56148 19616 56160
rect 19392 56120 19616 56148
rect 19392 56108 19398 56120
rect 19610 56108 19616 56120
rect 19668 56108 19674 56160
rect 19702 56108 19708 56160
rect 19760 56148 19766 56160
rect 19797 56151 19855 56157
rect 19797 56148 19809 56151
rect 19760 56120 19809 56148
rect 19760 56108 19766 56120
rect 19797 56117 19809 56120
rect 19843 56117 19855 56151
rect 19797 56111 19855 56117
rect 19886 56108 19892 56160
rect 19944 56108 19950 56160
rect 19996 56148 20024 56188
rect 22066 56160 22094 56188
rect 22557 56185 22569 56219
rect 22603 56185 22615 56219
rect 23308 56216 23336 56247
rect 24964 56216 24992 56247
rect 23308 56188 24992 56216
rect 25593 56219 25651 56225
rect 22557 56179 22615 56185
rect 25593 56185 25605 56219
rect 25639 56216 25651 56219
rect 25884 56216 25912 56299
rect 26160 56293 26188 56392
rect 27062 56380 27068 56392
rect 27120 56380 27126 56432
rect 27706 56420 27712 56432
rect 27264 56392 27712 56420
rect 26421 56355 26479 56361
rect 26421 56321 26433 56355
rect 26467 56321 26479 56355
rect 26421 56315 26479 56321
rect 26145 56287 26203 56293
rect 26145 56253 26157 56287
rect 26191 56253 26203 56287
rect 26436 56284 26464 56315
rect 27154 56312 27160 56364
rect 27212 56312 27218 56364
rect 27264 56284 27292 56392
rect 27706 56380 27712 56392
rect 27764 56380 27770 56432
rect 30098 56420 30104 56432
rect 27816 56392 30104 56420
rect 27816 56361 27844 56392
rect 30098 56380 30104 56392
rect 30156 56380 30162 56432
rect 27801 56355 27859 56361
rect 27801 56321 27813 56355
rect 27847 56321 27859 56355
rect 27801 56315 27859 56321
rect 28629 56355 28687 56361
rect 28629 56321 28641 56355
rect 28675 56352 28687 56355
rect 31757 56355 31815 56361
rect 28675 56324 31616 56352
rect 28675 56321 28687 56324
rect 28629 56315 28687 56321
rect 26436 56256 27292 56284
rect 27525 56287 27583 56293
rect 26145 56247 26203 56253
rect 27525 56253 27537 56287
rect 27571 56253 27583 56287
rect 27525 56247 27583 56253
rect 25639 56188 25912 56216
rect 26160 56216 26188 56247
rect 27540 56216 27568 56247
rect 28718 56244 28724 56296
rect 28776 56244 28782 56296
rect 28813 56287 28871 56293
rect 28813 56253 28825 56287
rect 28859 56253 28871 56287
rect 31588 56284 31616 56324
rect 31757 56321 31769 56355
rect 31803 56352 31815 56355
rect 32140 56352 32168 56451
rect 32214 56448 32220 56500
rect 32272 56488 32278 56500
rect 32490 56488 32496 56500
rect 32272 56460 32496 56488
rect 32272 56448 32278 56460
rect 32490 56448 32496 56460
rect 32548 56488 32554 56500
rect 32585 56491 32643 56497
rect 32585 56488 32597 56491
rect 32548 56460 32597 56488
rect 32548 56448 32554 56460
rect 32585 56457 32597 56460
rect 32631 56457 32643 56491
rect 32585 56451 32643 56457
rect 34701 56491 34759 56497
rect 34701 56457 34713 56491
rect 34747 56488 34759 56491
rect 35894 56488 35900 56500
rect 34747 56460 34928 56488
rect 34747 56457 34759 56460
rect 34701 56451 34759 56457
rect 31803 56324 32168 56352
rect 32493 56355 32551 56361
rect 31803 56321 31815 56324
rect 31757 56315 31815 56321
rect 32493 56321 32505 56355
rect 32539 56352 32551 56355
rect 34333 56355 34391 56361
rect 32539 56324 34284 56352
rect 32539 56321 32551 56324
rect 32493 56315 32551 56321
rect 34256 56296 34284 56324
rect 34333 56321 34345 56355
rect 34379 56321 34391 56355
rect 34900 56352 34928 56460
rect 35866 56448 35900 56488
rect 35952 56488 35958 56500
rect 36633 56491 36691 56497
rect 36633 56488 36645 56491
rect 35952 56460 36645 56488
rect 35952 56448 35958 56460
rect 36633 56457 36645 56460
rect 36679 56457 36691 56491
rect 38102 56488 38108 56500
rect 36633 56451 36691 56457
rect 36740 56460 38108 56488
rect 34977 56355 35035 56361
rect 34977 56352 34989 56355
rect 34900 56324 34989 56352
rect 34333 56315 34391 56321
rect 34977 56321 34989 56324
rect 35023 56321 35035 56355
rect 35866 56352 35894 56448
rect 34977 56315 35035 56321
rect 35084 56324 35894 56352
rect 32214 56284 32220 56296
rect 31588 56256 32220 56284
rect 28813 56247 28871 56253
rect 28828 56216 28856 56247
rect 32214 56244 32220 56256
rect 32272 56244 32278 56296
rect 32674 56244 32680 56296
rect 32732 56284 32738 56296
rect 34057 56287 34115 56293
rect 34057 56284 34069 56287
rect 32732 56256 34069 56284
rect 32732 56244 32738 56256
rect 34057 56253 34069 56256
rect 34103 56253 34115 56287
rect 34057 56247 34115 56253
rect 26160 56188 28856 56216
rect 34072 56216 34100 56247
rect 34238 56244 34244 56296
rect 34296 56244 34302 56296
rect 34348 56284 34376 56315
rect 35084 56284 35112 56324
rect 36262 56312 36268 56364
rect 36320 56352 36326 56364
rect 36740 56361 36768 56460
rect 38102 56448 38108 56460
rect 38160 56488 38166 56500
rect 38381 56491 38439 56497
rect 38381 56488 38393 56491
rect 38160 56460 38393 56488
rect 38160 56448 38166 56460
rect 38381 56457 38393 56460
rect 38427 56457 38439 56491
rect 38381 56451 38439 56457
rect 38473 56491 38531 56497
rect 38473 56457 38485 56491
rect 38519 56488 38531 56491
rect 40218 56488 40224 56500
rect 38519 56460 40224 56488
rect 38519 56457 38531 56460
rect 38473 56451 38531 56457
rect 40218 56448 40224 56460
rect 40276 56488 40282 56500
rect 40313 56491 40371 56497
rect 40313 56488 40325 56491
rect 40276 56460 40325 56488
rect 40276 56448 40282 56460
rect 40313 56457 40325 56460
rect 40359 56457 40371 56491
rect 40313 56451 40371 56457
rect 42429 56491 42487 56497
rect 42429 56457 42441 56491
rect 42475 56457 42487 56491
rect 42429 56451 42487 56457
rect 49237 56491 49295 56497
rect 49237 56457 49249 56491
rect 49283 56488 49295 56491
rect 49418 56488 49424 56500
rect 49283 56460 49424 56488
rect 49283 56457 49295 56460
rect 49237 56451 49295 56457
rect 37016 56392 40172 56420
rect 36725 56355 36783 56361
rect 36725 56352 36737 56355
rect 36320 56324 36737 56352
rect 36320 56312 36326 56324
rect 36725 56321 36737 56324
rect 36771 56321 36783 56355
rect 36725 56315 36783 56321
rect 36449 56287 36507 56293
rect 36449 56284 36461 56287
rect 34348 56256 35112 56284
rect 35866 56256 36461 56284
rect 35866 56216 35894 56256
rect 36449 56253 36461 56256
rect 36495 56284 36507 56287
rect 37016 56284 37044 56392
rect 37277 56355 37335 56361
rect 37277 56352 37289 56355
rect 36495 56256 37044 56284
rect 37200 56324 37289 56352
rect 36495 56253 36507 56256
rect 36449 56247 36507 56253
rect 34072 56188 35894 56216
rect 37093 56219 37151 56225
rect 25639 56185 25651 56188
rect 25593 56179 25651 56185
rect 37093 56185 37105 56219
rect 37139 56216 37151 56219
rect 37200 56216 37228 56324
rect 37277 56321 37289 56324
rect 37323 56321 37335 56355
rect 37277 56315 37335 56321
rect 38212 56293 38240 56392
rect 39117 56355 39175 56361
rect 39117 56352 39129 56355
rect 38856 56324 39129 56352
rect 38197 56287 38255 56293
rect 38197 56253 38209 56287
rect 38243 56253 38255 56287
rect 38197 56247 38255 56253
rect 38856 56225 38884 56324
rect 39117 56321 39129 56324
rect 39163 56321 39175 56355
rect 39117 56315 39175 56321
rect 39577 56355 39635 56361
rect 39577 56321 39589 56355
rect 39623 56352 39635 56355
rect 39623 56324 39896 56352
rect 39623 56321 39635 56324
rect 39577 56315 39635 56321
rect 39868 56225 39896 56324
rect 40144 56284 40172 56392
rect 40221 56355 40279 56361
rect 40221 56321 40233 56355
rect 40267 56352 40279 56355
rect 41509 56355 41567 56361
rect 40267 56324 41460 56352
rect 40267 56321 40279 56324
rect 40221 56315 40279 56321
rect 40405 56287 40463 56293
rect 40405 56284 40417 56287
rect 40144 56256 40417 56284
rect 40405 56253 40417 56256
rect 40451 56253 40463 56287
rect 41432 56284 41460 56324
rect 41509 56321 41521 56355
rect 41555 56352 41567 56355
rect 42444 56352 42472 56451
rect 42797 56423 42855 56429
rect 42797 56389 42809 56423
rect 42843 56420 42855 56423
rect 43898 56420 43904 56432
rect 42843 56392 43904 56420
rect 42843 56389 42855 56392
rect 42797 56383 42855 56389
rect 43898 56380 43904 56392
rect 43956 56380 43962 56432
rect 44453 56423 44511 56429
rect 44453 56389 44465 56423
rect 44499 56420 44511 56423
rect 45373 56423 45431 56429
rect 45373 56420 45385 56423
rect 44499 56392 45385 56420
rect 44499 56389 44511 56392
rect 44453 56383 44511 56389
rect 45373 56389 45385 56392
rect 45419 56420 45431 56423
rect 46934 56420 46940 56432
rect 45419 56392 46940 56420
rect 45419 56389 45431 56392
rect 45373 56383 45431 56389
rect 46934 56380 46940 56392
rect 46992 56420 46998 56432
rect 47670 56420 47676 56432
rect 46992 56392 47676 56420
rect 46992 56380 46998 56392
rect 47670 56380 47676 56392
rect 47728 56380 47734 56432
rect 41555 56324 42472 56352
rect 43625 56355 43683 56361
rect 41555 56321 41567 56324
rect 41509 56315 41567 56321
rect 43625 56321 43637 56355
rect 43671 56352 43683 56355
rect 45281 56355 45339 56361
rect 43671 56324 44404 56352
rect 43671 56321 43683 56324
rect 43625 56315 43683 56321
rect 41598 56284 41604 56296
rect 41432 56256 41604 56284
rect 40405 56247 40463 56253
rect 37139 56188 37228 56216
rect 38841 56219 38899 56225
rect 37139 56185 37151 56188
rect 37093 56179 37151 56185
rect 38841 56185 38853 56219
rect 38887 56185 38899 56219
rect 38841 56179 38899 56185
rect 39853 56219 39911 56225
rect 39853 56185 39865 56219
rect 39899 56185 39911 56219
rect 40420 56216 40448 56247
rect 41598 56244 41604 56256
rect 41656 56284 41662 56296
rect 41966 56284 41972 56296
rect 41656 56256 41972 56284
rect 41656 56244 41662 56256
rect 41966 56244 41972 56256
rect 42024 56284 42030 56296
rect 42889 56287 42947 56293
rect 42889 56284 42901 56287
rect 42024 56256 42901 56284
rect 42024 56244 42030 56256
rect 42889 56253 42901 56256
rect 42935 56253 42947 56287
rect 42889 56247 42947 56253
rect 42981 56287 43039 56293
rect 42981 56253 42993 56287
rect 43027 56253 43039 56287
rect 42981 56247 43039 56253
rect 42996 56216 43024 56247
rect 43714 56244 43720 56296
rect 43772 56244 43778 56296
rect 44376 56293 44404 56324
rect 45281 56321 45293 56355
rect 45327 56352 45339 56355
rect 45830 56352 45836 56364
rect 45327 56324 45836 56352
rect 45327 56321 45339 56324
rect 45281 56315 45339 56321
rect 45830 56312 45836 56324
rect 45888 56352 45894 56364
rect 49252 56352 49280 56451
rect 49418 56448 49424 56460
rect 49476 56448 49482 56500
rect 49786 56448 49792 56500
rect 49844 56448 49850 56500
rect 51445 56491 51503 56497
rect 51445 56457 51457 56491
rect 51491 56488 51503 56491
rect 51994 56488 52000 56500
rect 51491 56460 52000 56488
rect 51491 56457 51503 56460
rect 51445 56451 51503 56457
rect 51994 56448 52000 56460
rect 52052 56488 52058 56500
rect 52546 56488 52552 56500
rect 52052 56460 52552 56488
rect 52052 56448 52058 56460
rect 52546 56448 52552 56460
rect 52604 56448 52610 56500
rect 52730 56448 52736 56500
rect 52788 56448 52794 56500
rect 49329 56423 49387 56429
rect 49329 56389 49341 56423
rect 49375 56389 49387 56423
rect 51166 56420 51172 56432
rect 49329 56383 49387 56389
rect 49896 56392 51172 56420
rect 45888 56324 49280 56352
rect 49344 56352 49372 56383
rect 49896 56352 49924 56392
rect 51166 56380 51172 56392
rect 51224 56420 51230 56432
rect 51353 56423 51411 56429
rect 51353 56420 51365 56423
rect 51224 56392 51365 56420
rect 51224 56380 51230 56392
rect 51353 56389 51365 56392
rect 51399 56389 51411 56423
rect 51353 56383 51411 56389
rect 52914 56380 52920 56432
rect 52972 56420 52978 56432
rect 53193 56423 53251 56429
rect 53193 56420 53205 56423
rect 52972 56392 53205 56420
rect 52972 56380 52978 56392
rect 53193 56389 53205 56392
rect 53239 56420 53251 56423
rect 55214 56420 55220 56432
rect 53239 56392 55220 56420
rect 53239 56389 53251 56392
rect 53193 56383 53251 56389
rect 55214 56380 55220 56392
rect 55272 56420 55278 56432
rect 55858 56420 55864 56432
rect 55272 56392 55864 56420
rect 55272 56380 55278 56392
rect 55858 56380 55864 56392
rect 55916 56380 55922 56432
rect 49344 56324 49924 56352
rect 49973 56355 50031 56361
rect 45888 56312 45894 56324
rect 49973 56321 49985 56355
rect 50019 56321 50031 56355
rect 49973 56315 50031 56321
rect 50801 56355 50859 56361
rect 50801 56321 50813 56355
rect 50847 56352 50859 56355
rect 51074 56352 51080 56364
rect 50847 56324 51080 56352
rect 50847 56321 50859 56324
rect 50801 56315 50859 56321
rect 43809 56287 43867 56293
rect 43809 56253 43821 56287
rect 43855 56284 43867 56287
rect 44177 56287 44235 56293
rect 44177 56284 44189 56287
rect 43855 56256 44189 56284
rect 43855 56253 43867 56256
rect 43809 56247 43867 56253
rect 44177 56253 44189 56256
rect 44223 56253 44235 56287
rect 44177 56247 44235 56253
rect 44361 56287 44419 56293
rect 44361 56253 44373 56287
rect 44407 56284 44419 56287
rect 45002 56284 45008 56296
rect 44407 56256 45008 56284
rect 44407 56253 44419 56256
rect 44361 56247 44419 56253
rect 43824 56216 43852 56247
rect 40420 56188 43852 56216
rect 44192 56216 44220 56247
rect 45002 56244 45008 56256
rect 45060 56244 45066 56296
rect 45465 56287 45523 56293
rect 45465 56253 45477 56287
rect 45511 56253 45523 56287
rect 45465 56247 45523 56253
rect 45480 56216 45508 56247
rect 49050 56244 49056 56296
rect 49108 56244 49114 56296
rect 44192 56188 45508 56216
rect 49697 56219 49755 56225
rect 39853 56179 39911 56185
rect 49697 56185 49709 56219
rect 49743 56216 49755 56219
rect 49988 56216 50016 56315
rect 51074 56312 51080 56324
rect 51132 56312 51138 56364
rect 52089 56355 52147 56361
rect 52089 56352 52101 56355
rect 51828 56324 52101 56352
rect 51169 56287 51227 56293
rect 51169 56284 51181 56287
rect 49743 56188 50016 56216
rect 50632 56256 51181 56284
rect 49743 56185 49755 56188
rect 49697 56179 49755 56185
rect 20714 56148 20720 56160
rect 19996 56120 20720 56148
rect 20714 56108 20720 56120
rect 20772 56148 20778 56160
rect 21818 56148 21824 56160
rect 20772 56120 21824 56148
rect 20772 56108 20778 56120
rect 21818 56108 21824 56120
rect 21876 56108 21882 56160
rect 22066 56120 22100 56160
rect 22094 56108 22100 56120
rect 22152 56108 22158 56160
rect 22370 56108 22376 56160
rect 22428 56148 22434 56160
rect 22649 56151 22707 56157
rect 22649 56148 22661 56151
rect 22428 56120 22661 56148
rect 22428 56108 22434 56120
rect 22649 56117 22661 56120
rect 22695 56117 22707 56151
rect 22649 56111 22707 56117
rect 22738 56108 22744 56160
rect 22796 56148 22802 56160
rect 24029 56151 24087 56157
rect 24029 56148 24041 56151
rect 22796 56120 24041 56148
rect 22796 56108 22802 56120
rect 24029 56117 24041 56120
rect 24075 56117 24087 56151
rect 24029 56111 24087 56117
rect 25038 56108 25044 56160
rect 25096 56148 25102 56160
rect 25685 56151 25743 56157
rect 25685 56148 25697 56151
rect 25096 56120 25697 56148
rect 25096 56108 25102 56120
rect 25685 56117 25697 56120
rect 25731 56117 25743 56151
rect 25685 56111 25743 56117
rect 26970 56108 26976 56160
rect 27028 56108 27034 56160
rect 28074 56108 28080 56160
rect 28132 56148 28138 56160
rect 28261 56151 28319 56157
rect 28261 56148 28273 56151
rect 28132 56120 28273 56148
rect 28132 56108 28138 56120
rect 28261 56117 28273 56120
rect 28307 56117 28319 56151
rect 28261 56111 28319 56117
rect 31941 56151 31999 56157
rect 31941 56117 31953 56151
rect 31987 56148 31999 56151
rect 32398 56148 32404 56160
rect 31987 56120 32404 56148
rect 31987 56117 31999 56120
rect 31941 56111 31999 56117
rect 32398 56108 32404 56120
rect 32456 56108 32462 56160
rect 34790 56108 34796 56160
rect 34848 56108 34854 56160
rect 37461 56151 37519 56157
rect 37461 56117 37473 56151
rect 37507 56148 37519 56151
rect 37734 56148 37740 56160
rect 37507 56120 37740 56148
rect 37507 56117 37519 56120
rect 37461 56111 37519 56117
rect 37734 56108 37740 56120
rect 37792 56108 37798 56160
rect 38654 56108 38660 56160
rect 38712 56148 38718 56160
rect 38933 56151 38991 56157
rect 38933 56148 38945 56151
rect 38712 56120 38945 56148
rect 38712 56108 38718 56120
rect 38933 56117 38945 56120
rect 38979 56117 38991 56151
rect 38933 56111 38991 56117
rect 39761 56151 39819 56157
rect 39761 56117 39773 56151
rect 39807 56148 39819 56151
rect 40126 56148 40132 56160
rect 39807 56120 40132 56148
rect 39807 56117 39819 56120
rect 39761 56111 39819 56117
rect 40126 56108 40132 56120
rect 40184 56108 40190 56160
rect 41693 56151 41751 56157
rect 41693 56117 41705 56151
rect 41739 56148 41751 56151
rect 41966 56148 41972 56160
rect 41739 56120 41972 56148
rect 41739 56117 41751 56120
rect 41693 56111 41751 56117
rect 41966 56108 41972 56120
rect 42024 56108 42030 56160
rect 43257 56151 43315 56157
rect 43257 56117 43269 56151
rect 43303 56148 43315 56151
rect 43438 56148 43444 56160
rect 43303 56120 43444 56148
rect 43303 56117 43315 56120
rect 43257 56111 43315 56117
rect 43438 56108 43444 56120
rect 43496 56108 43502 56160
rect 44358 56108 44364 56160
rect 44416 56148 44422 56160
rect 44821 56151 44879 56157
rect 44821 56148 44833 56151
rect 44416 56120 44833 56148
rect 44416 56108 44422 56120
rect 44821 56117 44833 56120
rect 44867 56117 44879 56151
rect 44821 56111 44879 56117
rect 44910 56108 44916 56160
rect 44968 56108 44974 56160
rect 49050 56108 49056 56160
rect 49108 56148 49114 56160
rect 50632 56148 50660 56256
rect 51169 56253 51181 56256
rect 51215 56284 51227 56287
rect 51534 56284 51540 56296
rect 51215 56256 51540 56284
rect 51215 56253 51227 56256
rect 51169 56247 51227 56253
rect 51534 56244 51540 56256
rect 51592 56244 51598 56296
rect 50985 56219 51043 56225
rect 50985 56185 50997 56219
rect 51031 56216 51043 56219
rect 51718 56216 51724 56228
rect 51031 56188 51724 56216
rect 51031 56185 51043 56188
rect 50985 56179 51043 56185
rect 51718 56176 51724 56188
rect 51776 56176 51782 56228
rect 51828 56225 51856 56324
rect 52089 56321 52101 56324
rect 52135 56321 52147 56355
rect 52089 56315 52147 56321
rect 52365 56355 52423 56361
rect 52365 56321 52377 56355
rect 52411 56352 52423 56355
rect 52454 56352 52460 56364
rect 52411 56324 52460 56352
rect 52411 56321 52423 56324
rect 52365 56315 52423 56321
rect 52454 56312 52460 56324
rect 52512 56312 52518 56364
rect 53101 56355 53159 56361
rect 53101 56321 53113 56355
rect 53147 56352 53159 56355
rect 53561 56355 53619 56361
rect 53561 56352 53573 56355
rect 53147 56324 53573 56352
rect 53147 56321 53159 56324
rect 53101 56315 53159 56321
rect 53561 56321 53573 56324
rect 53607 56321 53619 56355
rect 53561 56315 53619 56321
rect 54205 56355 54263 56361
rect 54205 56321 54217 56355
rect 54251 56352 54263 56355
rect 55306 56352 55312 56364
rect 54251 56324 55312 56352
rect 54251 56321 54263 56324
rect 54205 56315 54263 56321
rect 55306 56312 55312 56324
rect 55364 56352 55370 56364
rect 56134 56352 56140 56364
rect 55364 56324 56140 56352
rect 55364 56312 55370 56324
rect 56134 56312 56140 56324
rect 56192 56312 56198 56364
rect 52270 56244 52276 56296
rect 52328 56284 52334 56296
rect 53285 56287 53343 56293
rect 53285 56284 53297 56287
rect 52328 56256 53297 56284
rect 52328 56244 52334 56256
rect 53285 56253 53297 56256
rect 53331 56253 53343 56287
rect 53285 56247 53343 56253
rect 51813 56219 51871 56225
rect 51813 56185 51825 56219
rect 51859 56185 51871 56219
rect 51813 56179 51871 56185
rect 49108 56120 50660 56148
rect 49108 56108 49114 56120
rect 51074 56108 51080 56160
rect 51132 56148 51138 56160
rect 51905 56151 51963 56157
rect 51905 56148 51917 56151
rect 51132 56120 51917 56148
rect 51132 56108 51138 56120
rect 51905 56117 51917 56120
rect 51951 56117 51963 56151
rect 51905 56111 51963 56117
rect 51994 56108 52000 56160
rect 52052 56148 52058 56160
rect 52181 56151 52239 56157
rect 52181 56148 52193 56151
rect 52052 56120 52193 56148
rect 52052 56108 52058 56120
rect 52181 56117 52193 56120
rect 52227 56117 52239 56151
rect 52181 56111 52239 56117
rect 1104 56058 58880 56080
rect 1104 56006 2350 56058
rect 2402 56006 2414 56058
rect 2466 56006 2478 56058
rect 2530 56006 2542 56058
rect 2594 56006 2606 56058
rect 2658 56006 33070 56058
rect 33122 56006 33134 56058
rect 33186 56006 33198 56058
rect 33250 56006 33262 56058
rect 33314 56006 33326 56058
rect 33378 56006 58880 56058
rect 1104 55984 58880 56006
rect 16577 55947 16635 55953
rect 16577 55913 16589 55947
rect 16623 55944 16635 55947
rect 16666 55944 16672 55956
rect 16623 55916 16672 55944
rect 16623 55913 16635 55916
rect 16577 55907 16635 55913
rect 16666 55904 16672 55916
rect 16724 55904 16730 55956
rect 18138 55904 18144 55956
rect 18196 55904 18202 55956
rect 18690 55904 18696 55956
rect 18748 55944 18754 55956
rect 19794 55944 19800 55956
rect 18748 55916 19800 55944
rect 18748 55904 18754 55916
rect 19794 55904 19800 55916
rect 19852 55904 19858 55956
rect 20888 55947 20946 55953
rect 20888 55913 20900 55947
rect 20934 55944 20946 55947
rect 22370 55944 22376 55956
rect 20934 55916 22376 55944
rect 20934 55913 20946 55916
rect 20888 55907 20946 55913
rect 22370 55904 22376 55916
rect 22428 55904 22434 55956
rect 43625 55947 43683 55953
rect 22572 55916 31754 55944
rect 16209 55879 16267 55885
rect 16209 55845 16221 55879
rect 16255 55876 16267 55879
rect 17862 55876 17868 55888
rect 16255 55848 17868 55876
rect 16255 55845 16267 55848
rect 16209 55839 16267 55845
rect 17862 55836 17868 55848
rect 17920 55836 17926 55888
rect 18509 55879 18567 55885
rect 18509 55845 18521 55879
rect 18555 55876 18567 55879
rect 19334 55876 19340 55888
rect 18555 55848 19340 55876
rect 18555 55845 18567 55848
rect 18509 55839 18567 55845
rect 19334 55836 19340 55848
rect 19392 55836 19398 55888
rect 19610 55836 19616 55888
rect 19668 55876 19674 55888
rect 20438 55876 20444 55888
rect 19668 55848 20444 55876
rect 19668 55836 19674 55848
rect 20438 55836 20444 55848
rect 20496 55836 20502 55888
rect 21910 55836 21916 55888
rect 21968 55876 21974 55888
rect 22572 55876 22600 55916
rect 21968 55848 22600 55876
rect 21968 55836 21974 55848
rect 23750 55836 23756 55888
rect 23808 55876 23814 55888
rect 24213 55879 24271 55885
rect 24213 55876 24225 55879
rect 23808 55848 24225 55876
rect 23808 55836 23814 55848
rect 24213 55845 24225 55848
rect 24259 55876 24271 55879
rect 24670 55876 24676 55888
rect 24259 55848 24676 55876
rect 24259 55845 24271 55848
rect 24213 55839 24271 55845
rect 24670 55836 24676 55848
rect 24728 55836 24734 55888
rect 27706 55836 27712 55888
rect 27764 55876 27770 55888
rect 27985 55879 28043 55885
rect 27985 55876 27997 55879
rect 27764 55848 27997 55876
rect 27764 55836 27770 55848
rect 27985 55845 27997 55848
rect 28031 55845 28043 55879
rect 27985 55839 28043 55845
rect 28718 55836 28724 55888
rect 28776 55876 28782 55888
rect 29549 55879 29607 55885
rect 29549 55876 29561 55879
rect 28776 55848 29561 55876
rect 28776 55836 28782 55848
rect 29549 55845 29561 55848
rect 29595 55845 29607 55879
rect 31726 55876 31754 55916
rect 43625 55913 43637 55947
rect 43671 55944 43683 55947
rect 43714 55944 43720 55956
rect 43671 55916 43720 55944
rect 43671 55913 43683 55916
rect 43625 55907 43683 55913
rect 43714 55904 43720 55916
rect 43772 55904 43778 55956
rect 45002 55904 45008 55956
rect 45060 55904 45066 55956
rect 52914 55944 52920 55956
rect 51276 55916 52920 55944
rect 32674 55876 32680 55888
rect 31726 55848 32680 55876
rect 29549 55839 29607 55845
rect 32674 55836 32680 55848
rect 32732 55836 32738 55888
rect 4062 55768 4068 55820
rect 4120 55808 4126 55820
rect 17129 55811 17187 55817
rect 4120 55780 17080 55808
rect 4120 55768 4126 55780
rect 15654 55700 15660 55752
rect 15712 55740 15718 55752
rect 15749 55743 15807 55749
rect 15749 55740 15761 55743
rect 15712 55712 15761 55740
rect 15712 55700 15718 55712
rect 15749 55709 15761 55712
rect 15795 55709 15807 55743
rect 15749 55703 15807 55709
rect 16022 55700 16028 55752
rect 16080 55700 16086 55752
rect 16301 55743 16359 55749
rect 16301 55709 16313 55743
rect 16347 55740 16359 55743
rect 16942 55740 16948 55752
rect 16347 55712 16948 55740
rect 16347 55709 16359 55712
rect 16301 55703 16359 55709
rect 16942 55700 16948 55712
rect 17000 55700 17006 55752
rect 17052 55740 17080 55780
rect 17129 55777 17141 55811
rect 17175 55808 17187 55811
rect 17310 55808 17316 55820
rect 17175 55780 17316 55808
rect 17175 55777 17187 55780
rect 17129 55771 17187 55777
rect 17310 55768 17316 55780
rect 17368 55768 17374 55820
rect 17586 55768 17592 55820
rect 17644 55768 17650 55820
rect 17681 55811 17739 55817
rect 17681 55777 17693 55811
rect 17727 55808 17739 55811
rect 18598 55808 18604 55820
rect 17727 55780 18604 55808
rect 17727 55777 17739 55780
rect 17681 55771 17739 55777
rect 17218 55740 17224 55752
rect 17052 55712 17224 55740
rect 17218 55700 17224 55712
rect 17276 55700 17282 55752
rect 16114 55632 16120 55684
rect 16172 55672 16178 55684
rect 17696 55672 17724 55771
rect 18598 55768 18604 55780
rect 18656 55768 18662 55820
rect 19518 55808 19524 55820
rect 19444 55780 19524 55808
rect 17770 55700 17776 55752
rect 17828 55700 17834 55752
rect 18322 55700 18328 55752
rect 18380 55700 18386 55752
rect 19444 55749 19472 55780
rect 19518 55768 19524 55780
rect 19576 55808 19582 55820
rect 20530 55808 20536 55820
rect 19576 55780 20536 55808
rect 19576 55768 19582 55780
rect 20530 55768 20536 55780
rect 20588 55768 20594 55820
rect 20625 55811 20683 55817
rect 20625 55777 20637 55811
rect 20671 55808 20683 55811
rect 22094 55808 22100 55820
rect 20671 55780 22100 55808
rect 20671 55777 20683 55780
rect 20625 55771 20683 55777
rect 22094 55768 22100 55780
rect 22152 55808 22158 55820
rect 22465 55811 22523 55817
rect 22465 55808 22477 55811
rect 22152 55780 22477 55808
rect 22152 55768 22158 55780
rect 22465 55777 22477 55780
rect 22511 55808 22523 55811
rect 24762 55808 24768 55820
rect 22511 55780 24768 55808
rect 22511 55777 22523 55780
rect 22465 55771 22523 55777
rect 24762 55768 24768 55780
rect 24820 55768 24826 55820
rect 26513 55811 26571 55817
rect 26513 55777 26525 55811
rect 26559 55808 26571 55811
rect 26970 55808 26976 55820
rect 26559 55780 26976 55808
rect 26559 55777 26571 55780
rect 26513 55771 26571 55777
rect 26970 55768 26976 55780
rect 27028 55768 27034 55820
rect 30098 55768 30104 55820
rect 30156 55768 30162 55820
rect 51276 55808 51304 55916
rect 52914 55904 52920 55916
rect 52972 55904 52978 55956
rect 53101 55947 53159 55953
rect 53101 55913 53113 55947
rect 53147 55944 53159 55947
rect 55306 55944 55312 55956
rect 53147 55916 55312 55944
rect 53147 55913 53159 55916
rect 53101 55907 53159 55913
rect 55306 55904 55312 55916
rect 55364 55904 55370 55956
rect 35866 55780 51304 55808
rect 18877 55743 18935 55749
rect 18877 55709 18889 55743
rect 18923 55740 18935 55743
rect 19245 55743 19303 55749
rect 19245 55740 19257 55743
rect 18923 55712 19257 55740
rect 18923 55709 18935 55712
rect 18877 55703 18935 55709
rect 19245 55709 19257 55712
rect 19291 55709 19303 55743
rect 19245 55703 19303 55709
rect 19429 55743 19487 55749
rect 19429 55709 19441 55743
rect 19475 55709 19487 55743
rect 19429 55703 19487 55709
rect 19702 55700 19708 55752
rect 19760 55700 19766 55752
rect 22002 55700 22008 55752
rect 22060 55700 22066 55752
rect 23842 55700 23848 55752
rect 23900 55740 23906 55752
rect 23900 55712 24808 55740
rect 23900 55700 23906 55712
rect 16172 55644 17724 55672
rect 16172 55632 16178 55644
rect 19610 55632 19616 55684
rect 19668 55632 19674 55684
rect 19812 55644 21312 55672
rect 15930 55564 15936 55616
rect 15988 55564 15994 55616
rect 16485 55607 16543 55613
rect 16485 55573 16497 55607
rect 16531 55604 16543 55607
rect 16758 55604 16764 55616
rect 16531 55576 16764 55604
rect 16531 55573 16543 55576
rect 16485 55567 16543 55573
rect 16758 55564 16764 55576
rect 16816 55564 16822 55616
rect 16942 55564 16948 55616
rect 17000 55564 17006 55616
rect 17037 55607 17095 55613
rect 17037 55573 17049 55607
rect 17083 55604 17095 55607
rect 17218 55604 17224 55616
rect 17083 55576 17224 55604
rect 17083 55573 17095 55576
rect 17037 55567 17095 55573
rect 17218 55564 17224 55576
rect 17276 55564 17282 55616
rect 19061 55607 19119 55613
rect 19061 55573 19073 55607
rect 19107 55604 19119 55607
rect 19812 55604 19840 55644
rect 19107 55576 19840 55604
rect 19889 55607 19947 55613
rect 19107 55573 19119 55576
rect 19061 55567 19119 55573
rect 19889 55573 19901 55607
rect 19935 55604 19947 55607
rect 20622 55604 20628 55616
rect 19935 55576 20628 55604
rect 19935 55573 19947 55576
rect 19889 55567 19947 55573
rect 20622 55564 20628 55576
rect 20680 55564 20686 55616
rect 21284 55604 21312 55644
rect 22296 55644 22508 55672
rect 22296 55604 22324 55644
rect 21284 55576 22324 55604
rect 22370 55564 22376 55616
rect 22428 55564 22434 55616
rect 22480 55604 22508 55644
rect 22738 55632 22744 55684
rect 22796 55632 22802 55684
rect 24780 55681 24808 55712
rect 26234 55700 26240 55752
rect 26292 55700 26298 55752
rect 28074 55700 28080 55752
rect 28132 55700 28138 55752
rect 35529 55743 35587 55749
rect 35529 55709 35541 55743
rect 35575 55740 35587 55743
rect 35866 55740 35894 55780
rect 35575 55712 35894 55740
rect 35575 55709 35587 55712
rect 35529 55703 35587 55709
rect 43438 55700 43444 55752
rect 43496 55700 43502 55752
rect 43898 55700 43904 55752
rect 43956 55740 43962 55752
rect 44177 55743 44235 55749
rect 44177 55740 44189 55743
rect 43956 55712 44189 55740
rect 43956 55700 43962 55712
rect 44177 55709 44189 55712
rect 44223 55709 44235 55743
rect 44177 55703 44235 55709
rect 44358 55700 44364 55752
rect 44416 55700 44422 55752
rect 44821 55743 44879 55749
rect 44821 55709 44833 55743
rect 44867 55740 44879 55743
rect 44910 55740 44916 55752
rect 44867 55712 44916 55740
rect 44867 55709 44879 55712
rect 44821 55703 44879 55709
rect 44910 55700 44916 55712
rect 44968 55700 44974 55752
rect 45554 55740 45560 55752
rect 45526 55700 45560 55740
rect 45612 55700 45618 55752
rect 24765 55675 24823 55681
rect 24044 55644 24532 55672
rect 23014 55604 23020 55616
rect 22480 55576 23020 55604
rect 23014 55564 23020 55576
rect 23072 55564 23078 55616
rect 23106 55564 23112 55616
rect 23164 55604 23170 55616
rect 24044 55604 24072 55644
rect 24504 55616 24532 55644
rect 24765 55641 24777 55675
rect 24811 55672 24823 55675
rect 26418 55672 26424 55684
rect 24811 55644 26424 55672
rect 24811 55641 24823 55644
rect 24765 55635 24823 55641
rect 26418 55632 26424 55644
rect 26476 55632 26482 55684
rect 27798 55672 27804 55684
rect 27738 55644 27804 55672
rect 27798 55632 27804 55644
rect 27856 55672 27862 55684
rect 27856 55644 29592 55672
rect 27856 55632 27862 55644
rect 29564 55616 29592 55644
rect 36170 55632 36176 55684
rect 36228 55672 36234 55684
rect 36265 55675 36323 55681
rect 36265 55672 36277 55675
rect 36228 55644 36277 55672
rect 36228 55632 36234 55644
rect 36265 55641 36277 55644
rect 36311 55641 36323 55675
rect 36265 55635 36323 55641
rect 38010 55632 38016 55684
rect 38068 55632 38074 55684
rect 44726 55632 44732 55684
rect 44784 55672 44790 55684
rect 45526 55672 45554 55700
rect 44784 55644 45554 55672
rect 51276 55672 51304 55780
rect 51626 55768 51632 55820
rect 51684 55768 51690 55820
rect 51350 55700 51356 55752
rect 51408 55700 51414 55752
rect 51276 55644 52118 55672
rect 44784 55632 44790 55644
rect 23164 55576 24072 55604
rect 23164 55564 23170 55576
rect 24486 55564 24492 55616
rect 24544 55564 24550 55616
rect 28261 55607 28319 55613
rect 28261 55573 28273 55607
rect 28307 55604 28319 55607
rect 28442 55604 28448 55616
rect 28307 55576 28448 55604
rect 28307 55573 28319 55576
rect 28261 55567 28319 55573
rect 28442 55564 28448 55576
rect 28500 55564 28506 55616
rect 29546 55564 29552 55616
rect 29604 55604 29610 55616
rect 33410 55604 33416 55616
rect 29604 55576 33416 55604
rect 29604 55564 29610 55576
rect 33410 55564 33416 55576
rect 33468 55604 33474 55616
rect 35437 55607 35495 55613
rect 35437 55604 35449 55607
rect 33468 55576 35449 55604
rect 33468 55564 33474 55576
rect 35437 55573 35449 55576
rect 35483 55604 35495 55607
rect 35526 55604 35532 55616
rect 35483 55576 35532 55604
rect 35483 55573 35495 55576
rect 35437 55567 35495 55573
rect 35526 55564 35532 55576
rect 35584 55564 35590 55616
rect 43254 55564 43260 55616
rect 43312 55564 43318 55616
rect 44542 55564 44548 55616
rect 44600 55564 44606 55616
rect 44634 55564 44640 55616
rect 44692 55564 44698 55616
rect 49602 55564 49608 55616
rect 49660 55604 49666 55616
rect 51534 55604 51540 55616
rect 49660 55576 51540 55604
rect 49660 55564 49666 55576
rect 51534 55564 51540 55576
rect 51592 55604 51598 55616
rect 52638 55604 52644 55616
rect 51592 55576 52644 55604
rect 51592 55564 51598 55576
rect 52638 55564 52644 55576
rect 52696 55564 52702 55616
rect 1104 55514 58880 55536
rect 1104 55462 3010 55514
rect 3062 55462 3074 55514
rect 3126 55462 3138 55514
rect 3190 55462 3202 55514
rect 3254 55462 3266 55514
rect 3318 55462 33730 55514
rect 33782 55462 33794 55514
rect 33846 55462 33858 55514
rect 33910 55462 33922 55514
rect 33974 55462 33986 55514
rect 34038 55462 58880 55514
rect 1104 55440 58880 55462
rect 17681 55403 17739 55409
rect 17681 55369 17693 55403
rect 17727 55400 17739 55403
rect 19702 55400 19708 55412
rect 17727 55372 19708 55400
rect 17727 55369 17739 55372
rect 17681 55363 17739 55369
rect 19702 55360 19708 55372
rect 19760 55360 19766 55412
rect 19794 55360 19800 55412
rect 19852 55400 19858 55412
rect 19889 55403 19947 55409
rect 19889 55400 19901 55403
rect 19852 55372 19901 55400
rect 19852 55360 19858 55372
rect 19889 55369 19901 55372
rect 19935 55369 19947 55403
rect 22094 55400 22100 55412
rect 19889 55363 19947 55369
rect 20088 55372 22100 55400
rect 16850 55292 16856 55344
rect 16908 55332 16914 55344
rect 19610 55332 19616 55344
rect 16908 55304 17172 55332
rect 19090 55304 19616 55332
rect 16908 55292 16914 55304
rect 16758 55224 16764 55276
rect 16816 55264 16822 55276
rect 17144 55273 17172 55304
rect 19610 55292 19616 55304
rect 19668 55292 19674 55344
rect 17129 55267 17187 55273
rect 16816 55236 17080 55264
rect 16816 55224 16822 55236
rect 16942 55156 16948 55208
rect 17000 55156 17006 55208
rect 17052 55128 17080 55236
rect 17129 55233 17141 55267
rect 17175 55233 17187 55267
rect 17129 55227 17187 55233
rect 17494 55224 17500 55276
rect 17552 55224 17558 55276
rect 19797 55267 19855 55273
rect 19797 55233 19809 55267
rect 19843 55264 19855 55267
rect 20088 55264 20116 55372
rect 22094 55360 22100 55372
rect 22152 55360 22158 55412
rect 22462 55360 22468 55412
rect 22520 55400 22526 55412
rect 26326 55400 26332 55412
rect 22520 55372 26332 55400
rect 22520 55360 22526 55372
rect 20898 55292 20904 55344
rect 20956 55332 20962 55344
rect 22002 55332 22008 55344
rect 20956 55304 22008 55332
rect 20956 55292 20962 55304
rect 22002 55292 22008 55304
rect 22060 55332 22066 55344
rect 23106 55332 23112 55344
rect 22060 55304 23112 55332
rect 22060 55292 22066 55304
rect 23106 55292 23112 55304
rect 23164 55292 23170 55344
rect 24486 55332 24492 55344
rect 23966 55304 24492 55332
rect 24486 55292 24492 55304
rect 24544 55292 24550 55344
rect 19843 55236 20116 55264
rect 21637 55267 21695 55273
rect 19843 55233 19855 55236
rect 19797 55227 19855 55233
rect 21637 55233 21649 55267
rect 21683 55264 21695 55267
rect 22094 55264 22100 55276
rect 21683 55236 22100 55264
rect 21683 55233 21695 55236
rect 21637 55227 21695 55233
rect 22094 55224 22100 55236
rect 22152 55224 22158 55276
rect 22278 55224 22284 55276
rect 22336 55264 22342 55276
rect 22465 55267 22523 55273
rect 22465 55264 22477 55267
rect 22336 55236 22477 55264
rect 22336 55224 22342 55236
rect 22465 55233 22477 55236
rect 22511 55233 22523 55267
rect 22465 55227 22523 55233
rect 22830 55224 22836 55276
rect 22888 55224 22894 55276
rect 23014 55224 23020 55276
rect 23072 55264 23078 55276
rect 24673 55267 24731 55273
rect 23072 55236 23244 55264
rect 23072 55224 23078 55236
rect 17954 55156 17960 55208
rect 18012 55196 18018 55208
rect 18049 55199 18107 55205
rect 18049 55196 18061 55199
rect 18012 55168 18061 55196
rect 18012 55156 18018 55168
rect 18049 55165 18061 55168
rect 18095 55165 18107 55199
rect 19521 55199 19579 55205
rect 19521 55196 19533 55199
rect 18049 55159 18107 55165
rect 18156 55168 19533 55196
rect 18156 55128 18184 55168
rect 19521 55165 19533 55168
rect 19567 55165 19579 55199
rect 19521 55159 19579 55165
rect 19886 55156 19892 55208
rect 19944 55196 19950 55208
rect 21361 55199 21419 55205
rect 21361 55196 21373 55199
rect 19944 55168 21373 55196
rect 19944 55156 19950 55168
rect 21361 55165 21373 55168
rect 21407 55165 21419 55199
rect 21361 55159 21419 55165
rect 21818 55156 21824 55208
rect 21876 55156 21882 55208
rect 22848 55196 22876 55224
rect 22925 55199 22983 55205
rect 22925 55196 22937 55199
rect 22848 55168 22937 55196
rect 22925 55165 22937 55168
rect 22971 55165 22983 55199
rect 23216 55196 23244 55236
rect 24673 55233 24685 55267
rect 24719 55264 24731 55267
rect 24780 55264 24808 55372
rect 26326 55360 26332 55372
rect 26384 55360 26390 55412
rect 26513 55403 26571 55409
rect 26513 55369 26525 55403
rect 26559 55400 26571 55403
rect 27062 55400 27068 55412
rect 26559 55372 27068 55400
rect 26559 55369 26571 55372
rect 26513 55363 26571 55369
rect 27062 55360 27068 55372
rect 27120 55360 27126 55412
rect 29917 55403 29975 55409
rect 28184 55372 29776 55400
rect 25038 55292 25044 55344
rect 25096 55292 25102 55344
rect 26418 55332 26424 55344
rect 26266 55304 26424 55332
rect 26418 55292 26424 55304
rect 26476 55332 26482 55344
rect 27798 55332 27804 55344
rect 26476 55304 27804 55332
rect 26476 55292 26482 55304
rect 27798 55292 27804 55304
rect 27856 55292 27862 55344
rect 26510 55264 26516 55276
rect 24719 55236 24808 55264
rect 26252 55236 26516 55264
rect 24719 55233 24731 55236
rect 24673 55227 24731 55233
rect 24397 55199 24455 55205
rect 24397 55196 24409 55199
rect 23216 55168 24409 55196
rect 22925 55159 22983 55165
rect 24397 55165 24409 55168
rect 24443 55165 24455 55199
rect 24397 55159 24455 55165
rect 24762 55156 24768 55208
rect 24820 55156 24826 55208
rect 17052 55100 18184 55128
rect 19978 55020 19984 55072
rect 20036 55060 20042 55072
rect 23290 55060 23296 55072
rect 20036 55032 23296 55060
rect 20036 55020 20042 55032
rect 23290 55020 23296 55032
rect 23348 55020 23354 55072
rect 24780 55060 24808 55156
rect 26252 55060 26280 55236
rect 26510 55224 26516 55236
rect 26568 55264 26574 55276
rect 28184 55273 28212 55372
rect 28442 55292 28448 55344
rect 28500 55292 28506 55344
rect 28169 55267 28227 55273
rect 28169 55264 28181 55267
rect 26568 55236 28181 55264
rect 26568 55224 26574 55236
rect 28169 55233 28181 55236
rect 28215 55233 28227 55267
rect 28169 55227 28227 55233
rect 29546 55224 29552 55276
rect 29604 55224 29610 55276
rect 29748 55264 29776 55372
rect 29917 55369 29929 55403
rect 29963 55400 29975 55403
rect 32030 55400 32036 55412
rect 29963 55372 32036 55400
rect 29963 55369 29975 55372
rect 29917 55363 29975 55369
rect 32030 55360 32036 55372
rect 32088 55360 32094 55412
rect 35713 55403 35771 55409
rect 32140 55372 33824 55400
rect 32140 55273 32168 55372
rect 32398 55292 32404 55344
rect 32456 55292 32462 55344
rect 33410 55292 33416 55344
rect 33468 55292 33474 55344
rect 32125 55267 32183 55273
rect 32125 55264 32137 55267
rect 29748 55236 32137 55264
rect 32125 55233 32137 55236
rect 32171 55233 32183 55267
rect 33796 55264 33824 55372
rect 35713 55369 35725 55403
rect 35759 55400 35771 55403
rect 35894 55400 35900 55412
rect 35759 55372 35900 55400
rect 35759 55369 35771 55372
rect 35713 55363 35771 55369
rect 35894 55360 35900 55372
rect 35952 55360 35958 55412
rect 37918 55360 37924 55412
rect 37976 55400 37982 55412
rect 38470 55400 38476 55412
rect 37976 55372 38476 55400
rect 37976 55360 37982 55372
rect 38470 55360 38476 55372
rect 38528 55360 38534 55412
rect 39761 55403 39819 55409
rect 38672 55372 39712 55400
rect 35526 55332 35532 55344
rect 35466 55304 35532 55332
rect 35526 55292 35532 55304
rect 35584 55292 35590 55344
rect 37274 55292 37280 55344
rect 37332 55332 37338 55344
rect 38672 55332 38700 55372
rect 39684 55332 39712 55372
rect 39761 55369 39773 55403
rect 39807 55400 39819 55403
rect 40218 55400 40224 55412
rect 39807 55372 40224 55400
rect 39807 55369 39819 55372
rect 39761 55363 39819 55369
rect 40218 55360 40224 55372
rect 40276 55360 40282 55412
rect 40512 55372 41460 55400
rect 40512 55332 40540 55372
rect 41432 55332 41460 55372
rect 41598 55360 41604 55412
rect 41656 55360 41662 55412
rect 43180 55372 43392 55400
rect 43180 55332 43208 55372
rect 37332 55304 38778 55332
rect 39684 55304 40618 55332
rect 41432 55304 43208 55332
rect 37332 55292 37338 55304
rect 43254 55292 43260 55344
rect 43312 55292 43318 55344
rect 43364 55332 43392 55372
rect 43640 55372 44404 55400
rect 43640 55332 43668 55372
rect 43364 55304 43746 55332
rect 33965 55267 34023 55273
rect 33965 55264 33977 55267
rect 33796 55236 33977 55264
rect 32125 55227 32183 55233
rect 33965 55233 33977 55236
rect 34011 55233 34023 55267
rect 33965 55227 34023 55233
rect 37918 55224 37924 55276
rect 37976 55264 37982 55276
rect 39853 55267 39911 55273
rect 37976 55236 38056 55264
rect 37976 55224 37982 55236
rect 34241 55199 34299 55205
rect 34241 55165 34253 55199
rect 34287 55196 34299 55199
rect 34790 55196 34796 55208
rect 34287 55168 34796 55196
rect 34287 55165 34299 55168
rect 34241 55159 34299 55165
rect 34790 55156 34796 55168
rect 34848 55156 34854 55208
rect 38028 55205 38056 55236
rect 39853 55233 39865 55267
rect 39899 55233 39911 55267
rect 39853 55227 39911 55233
rect 38013 55199 38071 55205
rect 38013 55196 38025 55199
rect 37936 55168 38025 55196
rect 24780 55032 26280 55060
rect 33873 55063 33931 55069
rect 33873 55029 33885 55063
rect 33919 55060 33931 55063
rect 34238 55060 34244 55072
rect 33919 55032 34244 55060
rect 33919 55029 33931 55032
rect 33873 55023 33931 55029
rect 34238 55020 34244 55032
rect 34296 55020 34302 55072
rect 37936 55060 37964 55168
rect 38013 55165 38025 55168
rect 38059 55165 38071 55199
rect 38013 55159 38071 55165
rect 38378 55156 38384 55208
rect 38436 55196 38442 55208
rect 39868 55196 39896 55227
rect 38436 55168 39896 55196
rect 38436 55156 38442 55168
rect 39868 55140 39896 55168
rect 40126 55156 40132 55208
rect 40184 55156 40190 55208
rect 42978 55156 42984 55208
rect 43036 55156 43042 55208
rect 44266 55156 44272 55208
rect 44324 55196 44330 55208
rect 44376 55196 44404 55372
rect 44726 55360 44732 55412
rect 44784 55360 44790 55412
rect 46750 55400 46756 55412
rect 44836 55372 46756 55400
rect 44836 55273 44864 55372
rect 46750 55360 46756 55372
rect 46808 55360 46814 55412
rect 51350 55400 51356 55412
rect 48700 55372 51356 55400
rect 48590 55332 48596 55344
rect 46676 55304 48596 55332
rect 44821 55267 44879 55273
rect 44821 55233 44833 55267
rect 44867 55233 44879 55267
rect 46676 55264 46704 55304
rect 48590 55292 48596 55304
rect 48648 55292 48654 55344
rect 44821 55227 44879 55233
rect 46124 55236 46704 55264
rect 44324 55168 44404 55196
rect 44324 55156 44330 55168
rect 44542 55156 44548 55208
rect 44600 55196 44606 55208
rect 45097 55199 45155 55205
rect 45097 55196 45109 55199
rect 44600 55168 45109 55196
rect 44600 55156 44606 55168
rect 45097 55165 45109 55168
rect 45143 55165 45155 55199
rect 45097 55159 45155 55165
rect 45186 55156 45192 55208
rect 45244 55196 45250 55208
rect 46124 55196 46152 55236
rect 46750 55224 46756 55276
rect 46808 55264 46814 55276
rect 48700 55264 48728 55372
rect 48774 55292 48780 55344
rect 48832 55332 48838 55344
rect 49602 55332 49608 55344
rect 48832 55304 49608 55332
rect 48832 55292 48838 55304
rect 49602 55292 49608 55304
rect 49660 55292 49666 55344
rect 50816 55273 50844 55372
rect 51350 55360 51356 55372
rect 51408 55400 51414 55412
rect 54481 55403 54539 55409
rect 51408 55372 52776 55400
rect 51408 55360 51414 55372
rect 51074 55292 51080 55344
rect 51132 55292 51138 55344
rect 51534 55292 51540 55344
rect 51592 55292 51598 55344
rect 52748 55273 52776 55372
rect 54481 55369 54493 55403
rect 54527 55400 54539 55403
rect 55214 55400 55220 55412
rect 54527 55372 55220 55400
rect 54527 55369 54539 55372
rect 54481 55363 54539 55369
rect 55214 55360 55220 55372
rect 55272 55360 55278 55412
rect 52914 55292 52920 55344
rect 52972 55332 52978 55344
rect 53466 55332 53472 55344
rect 52972 55304 53472 55332
rect 52972 55292 52978 55304
rect 53466 55292 53472 55304
rect 53524 55292 53530 55344
rect 48869 55267 48927 55273
rect 48869 55264 48881 55267
rect 46808 55236 48881 55264
rect 46808 55224 46814 55236
rect 48869 55233 48881 55236
rect 48915 55233 48927 55267
rect 48869 55227 48927 55233
rect 50801 55267 50859 55273
rect 50801 55233 50813 55267
rect 50847 55233 50859 55267
rect 50801 55227 50859 55233
rect 52733 55267 52791 55273
rect 52733 55233 52745 55267
rect 52779 55233 52791 55267
rect 52733 55227 52791 55233
rect 45244 55168 46152 55196
rect 46569 55199 46627 55205
rect 45244 55156 45250 55168
rect 46569 55165 46581 55199
rect 46615 55196 46627 55199
rect 46934 55196 46940 55208
rect 46615 55168 46940 55196
rect 46615 55165 46627 55168
rect 46569 55159 46627 55165
rect 46934 55156 46940 55168
rect 46992 55156 46998 55208
rect 49145 55199 49203 55205
rect 49145 55165 49157 55199
rect 49191 55196 49203 55199
rect 49786 55196 49792 55208
rect 49191 55168 49792 55196
rect 49191 55165 49203 55168
rect 49145 55159 49203 55165
rect 49786 55156 49792 55168
rect 49844 55156 49850 55208
rect 50617 55199 50675 55205
rect 50617 55165 50629 55199
rect 50663 55196 50675 55199
rect 51166 55196 51172 55208
rect 50663 55168 51172 55196
rect 50663 55165 50675 55168
rect 50617 55159 50675 55165
rect 51166 55156 51172 55168
rect 51224 55156 51230 55208
rect 51718 55156 51724 55208
rect 51776 55196 51782 55208
rect 51776 55168 52132 55196
rect 51776 55156 51782 55168
rect 39850 55088 39856 55140
rect 39908 55088 39914 55140
rect 52104 55128 52132 55168
rect 52546 55156 52552 55208
rect 52604 55156 52610 55208
rect 53009 55199 53067 55205
rect 53009 55196 53021 55199
rect 52656 55168 53021 55196
rect 52656 55128 52684 55168
rect 53009 55165 53021 55168
rect 53055 55165 53067 55199
rect 53009 55159 53067 55165
rect 52104 55100 52684 55128
rect 38010 55060 38016 55072
rect 37936 55032 38016 55060
rect 38010 55020 38016 55032
rect 38068 55020 38074 55072
rect 38276 55063 38334 55069
rect 38276 55029 38288 55063
rect 38322 55060 38334 55063
rect 38654 55060 38660 55072
rect 38322 55032 38660 55060
rect 38322 55029 38334 55032
rect 38276 55023 38334 55029
rect 38654 55020 38660 55032
rect 38712 55020 38718 55072
rect 1104 54970 58880 54992
rect 1104 54918 2350 54970
rect 2402 54918 2414 54970
rect 2466 54918 2478 54970
rect 2530 54918 2542 54970
rect 2594 54918 2606 54970
rect 2658 54918 33070 54970
rect 33122 54918 33134 54970
rect 33186 54918 33198 54970
rect 33250 54918 33262 54970
rect 33314 54918 33326 54970
rect 33378 54918 58880 54970
rect 1104 54896 58880 54918
rect 20438 54816 20444 54868
rect 20496 54856 20502 54868
rect 20625 54859 20683 54865
rect 20625 54856 20637 54859
rect 20496 54828 20637 54856
rect 20496 54816 20502 54828
rect 20625 54825 20637 54828
rect 20671 54825 20683 54859
rect 20625 54819 20683 54825
rect 20732 54828 22600 54856
rect 19334 54748 19340 54800
rect 19392 54788 19398 54800
rect 20732 54788 20760 54828
rect 19392 54760 20760 54788
rect 19392 54748 19398 54760
rect 22373 54723 22431 54729
rect 22373 54689 22385 54723
rect 22419 54720 22431 54723
rect 22462 54720 22468 54732
rect 22419 54692 22468 54720
rect 22419 54689 22431 54692
rect 22373 54683 22431 54689
rect 22462 54680 22468 54692
rect 22520 54680 22526 54732
rect 22572 54720 22600 54828
rect 23290 54816 23296 54868
rect 23348 54856 23354 54868
rect 24213 54859 24271 54865
rect 24213 54856 24225 54859
rect 23348 54828 24225 54856
rect 23348 54816 23354 54828
rect 24213 54825 24225 54828
rect 24259 54825 24271 54859
rect 24213 54819 24271 54825
rect 29365 54859 29423 54865
rect 29365 54825 29377 54859
rect 29411 54856 29423 54859
rect 30098 54856 30104 54868
rect 29411 54828 30104 54856
rect 29411 54825 29423 54828
rect 29365 54819 29423 54825
rect 30098 54816 30104 54828
rect 30156 54816 30162 54868
rect 36262 54816 36268 54868
rect 36320 54816 36326 54868
rect 39850 54816 39856 54868
rect 39908 54856 39914 54868
rect 41141 54859 41199 54865
rect 41141 54856 41153 54859
rect 39908 54828 41153 54856
rect 39908 54816 39914 54828
rect 41141 54825 41153 54828
rect 41187 54825 41199 54859
rect 41141 54819 41199 54825
rect 43441 54859 43499 54865
rect 43441 54825 43453 54859
rect 43487 54856 43499 54859
rect 43898 54856 43904 54868
rect 43487 54828 43904 54856
rect 43487 54825 43499 54828
rect 43441 54819 43499 54825
rect 26234 54748 26240 54800
rect 26292 54748 26298 54800
rect 22741 54723 22799 54729
rect 22741 54720 22753 54723
rect 22572 54692 22753 54720
rect 22741 54689 22753 54692
rect 22787 54689 22799 54723
rect 26252 54720 26280 54748
rect 27617 54723 27675 54729
rect 27617 54720 27629 54723
rect 26252 54692 27629 54720
rect 22741 54683 22799 54689
rect 27617 54689 27629 54692
rect 27663 54689 27675 54723
rect 27617 54683 27675 54689
rect 27890 54680 27896 54732
rect 27948 54680 27954 54732
rect 37734 54680 37740 54732
rect 37792 54680 37798 54732
rect 38010 54680 38016 54732
rect 38068 54680 38074 54732
rect 41156 54720 41184 54819
rect 43898 54816 43904 54828
rect 43956 54816 43962 54868
rect 53006 54816 53012 54868
rect 53064 54856 53070 54868
rect 53101 54859 53159 54865
rect 53101 54856 53113 54859
rect 53064 54828 53113 54856
rect 53064 54816 53070 54828
rect 53101 54825 53113 54828
rect 53147 54825 53159 54859
rect 53101 54819 53159 54825
rect 41693 54723 41751 54729
rect 41693 54720 41705 54723
rect 41156 54692 41705 54720
rect 41693 54689 41705 54692
rect 41739 54720 41751 54723
rect 42978 54720 42984 54732
rect 41739 54692 42984 54720
rect 41739 54689 41751 54692
rect 41693 54683 41751 54689
rect 42978 54680 42984 54692
rect 43036 54680 43042 54732
rect 46750 54680 46756 54732
rect 46808 54680 46814 54732
rect 51350 54680 51356 54732
rect 51408 54680 51414 54732
rect 51629 54723 51687 54729
rect 51629 54689 51641 54723
rect 51675 54720 51687 54723
rect 51994 54720 52000 54732
rect 51675 54692 52000 54720
rect 51675 54689 51687 54692
rect 51629 54683 51687 54689
rect 51994 54680 52000 54692
rect 52052 54680 52058 54732
rect 52638 54680 52644 54732
rect 52696 54720 52702 54732
rect 52696 54692 52960 54720
rect 52696 54680 52702 54692
rect 23842 54612 23848 54664
rect 23900 54612 23906 54664
rect 29546 54652 29552 54664
rect 29026 54624 29552 54652
rect 29546 54612 29552 54624
rect 29604 54612 29610 54664
rect 44266 54652 44272 54664
rect 43102 54624 44272 54652
rect 44266 54612 44272 54624
rect 44324 54652 44330 54664
rect 44818 54652 44824 54664
rect 44324 54624 44824 54652
rect 44324 54612 44330 54624
rect 44818 54612 44824 54624
rect 44876 54652 44882 54664
rect 45186 54652 45192 54664
rect 44876 54624 45192 54652
rect 44876 54612 44882 54624
rect 45186 54612 45192 54624
rect 45244 54612 45250 54664
rect 22002 54584 22008 54596
rect 21666 54556 22008 54584
rect 22002 54544 22008 54556
rect 22060 54544 22066 54596
rect 22097 54587 22155 54593
rect 22097 54553 22109 54587
rect 22143 54553 22155 54587
rect 22097 54547 22155 54553
rect 27525 54587 27583 54593
rect 27525 54553 27537 54587
rect 27571 54553 27583 54587
rect 36170 54584 36176 54596
rect 27525 54547 27583 54553
rect 29196 54556 36176 54584
rect 15930 54476 15936 54528
rect 15988 54516 15994 54528
rect 22112 54516 22140 54547
rect 15988 54488 22140 54516
rect 27540 54516 27568 54547
rect 27798 54516 27804 54528
rect 27540 54488 27804 54516
rect 15988 54476 15994 54488
rect 27798 54476 27804 54488
rect 27856 54516 27862 54528
rect 29196 54516 29224 54556
rect 36170 54544 36176 54556
rect 36228 54584 36234 54596
rect 36228 54556 36492 54584
rect 36228 54544 36234 54556
rect 27856 54488 29224 54516
rect 36464 54516 36492 54556
rect 37274 54544 37280 54596
rect 37332 54544 37338 54596
rect 39853 54587 39911 54593
rect 39853 54553 39865 54587
rect 39899 54553 39911 54587
rect 39853 54547 39911 54553
rect 39868 54516 39896 54547
rect 41966 54544 41972 54596
rect 42024 54544 42030 54596
rect 45005 54587 45063 54593
rect 45005 54584 45017 54587
rect 43272 54556 45017 54584
rect 43272 54516 43300 54556
rect 45005 54553 45017 54556
rect 45051 54553 45063 54587
rect 52932 54584 52960 54692
rect 53466 54612 53472 54664
rect 53524 54652 53530 54664
rect 53561 54655 53619 54661
rect 53561 54652 53573 54655
rect 53524 54624 53573 54652
rect 53524 54612 53530 54624
rect 53561 54621 53573 54624
rect 53607 54652 53619 54655
rect 58250 54652 58256 54664
rect 53607 54624 58256 54652
rect 53607 54621 53619 54624
rect 53561 54615 53619 54621
rect 58250 54612 58256 54624
rect 58308 54612 58314 54664
rect 53193 54587 53251 54593
rect 53193 54584 53205 54587
rect 52854 54556 53205 54584
rect 45005 54547 45063 54553
rect 53193 54553 53205 54556
rect 53239 54553 53251 54587
rect 53193 54547 53251 54553
rect 36464 54488 43300 54516
rect 27856 54476 27862 54488
rect 1104 54426 58880 54448
rect 1104 54374 3010 54426
rect 3062 54374 3074 54426
rect 3126 54374 3138 54426
rect 3190 54374 3202 54426
rect 3254 54374 3266 54426
rect 3318 54374 33730 54426
rect 33782 54374 33794 54426
rect 33846 54374 33858 54426
rect 33910 54374 33922 54426
rect 33974 54374 33986 54426
rect 34038 54374 58880 54426
rect 1104 54352 58880 54374
rect 19610 54272 19616 54324
rect 19668 54312 19674 54324
rect 46750 54312 46756 54324
rect 19668 54284 21036 54312
rect 19668 54272 19674 54284
rect 21008 54244 21036 54284
rect 44100 54284 46756 54312
rect 21082 54244 21088 54256
rect 20930 54216 21088 54244
rect 21082 54204 21088 54216
rect 21140 54244 21146 54256
rect 22002 54244 22008 54256
rect 21140 54216 22008 54244
rect 21140 54204 21146 54216
rect 22002 54204 22008 54216
rect 22060 54204 22066 54256
rect 44100 54185 44128 54284
rect 46750 54272 46756 54284
rect 46808 54272 46814 54324
rect 44361 54247 44419 54253
rect 44361 54213 44373 54247
rect 44407 54244 44419 54247
rect 44634 54244 44640 54256
rect 44407 54216 44640 54244
rect 44407 54213 44419 54216
rect 44361 54207 44419 54213
rect 44634 54204 44640 54216
rect 44692 54204 44698 54256
rect 44818 54204 44824 54256
rect 44876 54204 44882 54256
rect 44085 54179 44143 54185
rect 44085 54145 44097 54179
rect 44131 54145 44143 54179
rect 44085 54139 44143 54145
rect 20806 54068 20812 54120
rect 20864 54108 20870 54120
rect 21361 54111 21419 54117
rect 21361 54108 21373 54111
rect 20864 54080 21373 54108
rect 20864 54068 20870 54080
rect 21361 54077 21373 54080
rect 21407 54077 21419 54111
rect 21361 54071 21419 54077
rect 21637 54111 21695 54117
rect 21637 54077 21649 54111
rect 21683 54108 21695 54111
rect 22462 54108 22468 54120
rect 21683 54080 22468 54108
rect 21683 54077 21695 54080
rect 21637 54071 21695 54077
rect 22462 54068 22468 54080
rect 22520 54068 22526 54120
rect 45830 54068 45836 54120
rect 45888 54068 45894 54120
rect 16206 53932 16212 53984
rect 16264 53972 16270 53984
rect 19889 53975 19947 53981
rect 19889 53972 19901 53975
rect 16264 53944 19901 53972
rect 16264 53932 16270 53944
rect 19889 53941 19901 53944
rect 19935 53941 19947 53975
rect 19889 53935 19947 53941
rect 1104 53882 58880 53904
rect 1104 53830 2350 53882
rect 2402 53830 2414 53882
rect 2466 53830 2478 53882
rect 2530 53830 2542 53882
rect 2594 53830 2606 53882
rect 2658 53830 33070 53882
rect 33122 53830 33134 53882
rect 33186 53830 33198 53882
rect 33250 53830 33262 53882
rect 33314 53830 33326 53882
rect 33378 53830 58880 53882
rect 1104 53808 58880 53830
rect 17770 53728 17776 53780
rect 17828 53768 17834 53780
rect 20717 53771 20775 53777
rect 20717 53768 20729 53771
rect 17828 53740 20729 53768
rect 17828 53728 17834 53740
rect 20717 53737 20729 53740
rect 20763 53737 20775 53771
rect 20717 53731 20775 53737
rect 26510 53728 26516 53780
rect 26568 53728 26574 53780
rect 22462 53592 22468 53644
rect 22520 53592 22526 53644
rect 21082 53524 21088 53576
rect 21140 53524 21146 53576
rect 27798 53524 27804 53576
rect 27856 53524 27862 53576
rect 22189 53499 22247 53505
rect 22189 53465 22201 53499
rect 22235 53496 22247 53499
rect 22554 53496 22560 53508
rect 22235 53468 22560 53496
rect 22235 53465 22247 53468
rect 22189 53459 22247 53465
rect 22554 53456 22560 53468
rect 22612 53456 22618 53508
rect 1104 53338 58880 53360
rect 1104 53286 3010 53338
rect 3062 53286 3074 53338
rect 3126 53286 3138 53338
rect 3190 53286 3202 53338
rect 3254 53286 3266 53338
rect 3318 53286 33730 53338
rect 33782 53286 33794 53338
rect 33846 53286 33858 53338
rect 33910 53286 33922 53338
rect 33974 53286 33986 53338
rect 34038 53286 58880 53338
rect 1104 53264 58880 53286
rect 19426 53184 19432 53236
rect 19484 53224 19490 53236
rect 19613 53227 19671 53233
rect 19613 53224 19625 53227
rect 19484 53196 19625 53224
rect 19484 53184 19490 53196
rect 19613 53193 19625 53196
rect 19659 53193 19671 53227
rect 19613 53187 19671 53193
rect 21082 53156 21088 53168
rect 20654 53128 21088 53156
rect 21082 53116 21088 53128
rect 21140 53116 21146 53168
rect 21361 53091 21419 53097
rect 21361 53057 21373 53091
rect 21407 53088 21419 53091
rect 22462 53088 22468 53100
rect 21407 53060 22468 53088
rect 21407 53057 21419 53060
rect 21361 53051 21419 53057
rect 22462 53048 22468 53060
rect 22520 53048 22526 53100
rect 20622 52980 20628 53032
rect 20680 53020 20686 53032
rect 21085 53023 21143 53029
rect 21085 53020 21097 53023
rect 20680 52992 21097 53020
rect 20680 52980 20686 52992
rect 21085 52989 21097 52992
rect 21131 52989 21143 53023
rect 21085 52983 21143 52989
rect 1104 52794 58880 52816
rect 1104 52742 2350 52794
rect 2402 52742 2414 52794
rect 2466 52742 2478 52794
rect 2530 52742 2542 52794
rect 2594 52742 2606 52794
rect 2658 52742 33070 52794
rect 33122 52742 33134 52794
rect 33186 52742 33198 52794
rect 33250 52742 33262 52794
rect 33314 52742 33326 52794
rect 33378 52742 58880 52794
rect 1104 52720 58880 52742
rect 1104 52250 58880 52272
rect 1104 52198 3010 52250
rect 3062 52198 3074 52250
rect 3126 52198 3138 52250
rect 3190 52198 3202 52250
rect 3254 52198 3266 52250
rect 3318 52198 33730 52250
rect 33782 52198 33794 52250
rect 33846 52198 33858 52250
rect 33910 52198 33922 52250
rect 33974 52198 33986 52250
rect 34038 52198 58880 52250
rect 1104 52176 58880 52198
rect 1104 51706 58880 51728
rect 1104 51654 2350 51706
rect 2402 51654 2414 51706
rect 2466 51654 2478 51706
rect 2530 51654 2542 51706
rect 2594 51654 2606 51706
rect 2658 51654 33070 51706
rect 33122 51654 33134 51706
rect 33186 51654 33198 51706
rect 33250 51654 33262 51706
rect 33314 51654 33326 51706
rect 33378 51654 58880 51706
rect 1104 51632 58880 51654
rect 1104 51162 58880 51184
rect 1104 51110 3010 51162
rect 3062 51110 3074 51162
rect 3126 51110 3138 51162
rect 3190 51110 3202 51162
rect 3254 51110 3266 51162
rect 3318 51110 33730 51162
rect 33782 51110 33794 51162
rect 33846 51110 33858 51162
rect 33910 51110 33922 51162
rect 33974 51110 33986 51162
rect 34038 51110 58880 51162
rect 1104 51088 58880 51110
rect 1104 50618 58880 50640
rect 1104 50566 2350 50618
rect 2402 50566 2414 50618
rect 2466 50566 2478 50618
rect 2530 50566 2542 50618
rect 2594 50566 2606 50618
rect 2658 50566 33070 50618
rect 33122 50566 33134 50618
rect 33186 50566 33198 50618
rect 33250 50566 33262 50618
rect 33314 50566 33326 50618
rect 33378 50566 58880 50618
rect 1104 50544 58880 50566
rect 1104 50074 58880 50096
rect 1104 50022 3010 50074
rect 3062 50022 3074 50074
rect 3126 50022 3138 50074
rect 3190 50022 3202 50074
rect 3254 50022 3266 50074
rect 3318 50022 33730 50074
rect 33782 50022 33794 50074
rect 33846 50022 33858 50074
rect 33910 50022 33922 50074
rect 33974 50022 33986 50074
rect 34038 50022 58880 50074
rect 1104 50000 58880 50022
rect 1104 49530 58880 49552
rect 1104 49478 2350 49530
rect 2402 49478 2414 49530
rect 2466 49478 2478 49530
rect 2530 49478 2542 49530
rect 2594 49478 2606 49530
rect 2658 49478 33070 49530
rect 33122 49478 33134 49530
rect 33186 49478 33198 49530
rect 33250 49478 33262 49530
rect 33314 49478 33326 49530
rect 33378 49478 58880 49530
rect 1104 49456 58880 49478
rect 1104 48986 58880 49008
rect 1104 48934 3010 48986
rect 3062 48934 3074 48986
rect 3126 48934 3138 48986
rect 3190 48934 3202 48986
rect 3254 48934 3266 48986
rect 3318 48934 33730 48986
rect 33782 48934 33794 48986
rect 33846 48934 33858 48986
rect 33910 48934 33922 48986
rect 33974 48934 33986 48986
rect 34038 48934 58880 48986
rect 1104 48912 58880 48934
rect 1104 48442 58880 48464
rect 1104 48390 2350 48442
rect 2402 48390 2414 48442
rect 2466 48390 2478 48442
rect 2530 48390 2542 48442
rect 2594 48390 2606 48442
rect 2658 48390 33070 48442
rect 33122 48390 33134 48442
rect 33186 48390 33198 48442
rect 33250 48390 33262 48442
rect 33314 48390 33326 48442
rect 33378 48390 58880 48442
rect 1104 48368 58880 48390
rect 1104 47898 58880 47920
rect 1104 47846 3010 47898
rect 3062 47846 3074 47898
rect 3126 47846 3138 47898
rect 3190 47846 3202 47898
rect 3254 47846 3266 47898
rect 3318 47846 33730 47898
rect 33782 47846 33794 47898
rect 33846 47846 33858 47898
rect 33910 47846 33922 47898
rect 33974 47846 33986 47898
rect 34038 47846 58880 47898
rect 1104 47824 58880 47846
rect 1104 47354 58880 47376
rect 1104 47302 2350 47354
rect 2402 47302 2414 47354
rect 2466 47302 2478 47354
rect 2530 47302 2542 47354
rect 2594 47302 2606 47354
rect 2658 47302 33070 47354
rect 33122 47302 33134 47354
rect 33186 47302 33198 47354
rect 33250 47302 33262 47354
rect 33314 47302 33326 47354
rect 33378 47302 58880 47354
rect 1104 47280 58880 47302
rect 1104 46810 58880 46832
rect 1104 46758 3010 46810
rect 3062 46758 3074 46810
rect 3126 46758 3138 46810
rect 3190 46758 3202 46810
rect 3254 46758 3266 46810
rect 3318 46758 33730 46810
rect 33782 46758 33794 46810
rect 33846 46758 33858 46810
rect 33910 46758 33922 46810
rect 33974 46758 33986 46810
rect 34038 46758 58880 46810
rect 1104 46736 58880 46758
rect 1104 46266 58880 46288
rect 1104 46214 2350 46266
rect 2402 46214 2414 46266
rect 2466 46214 2478 46266
rect 2530 46214 2542 46266
rect 2594 46214 2606 46266
rect 2658 46214 33070 46266
rect 33122 46214 33134 46266
rect 33186 46214 33198 46266
rect 33250 46214 33262 46266
rect 33314 46214 33326 46266
rect 33378 46214 58880 46266
rect 1104 46192 58880 46214
rect 1104 45722 58880 45744
rect 1104 45670 3010 45722
rect 3062 45670 3074 45722
rect 3126 45670 3138 45722
rect 3190 45670 3202 45722
rect 3254 45670 3266 45722
rect 3318 45670 33730 45722
rect 33782 45670 33794 45722
rect 33846 45670 33858 45722
rect 33910 45670 33922 45722
rect 33974 45670 33986 45722
rect 34038 45670 58880 45722
rect 1104 45648 58880 45670
rect 1104 45178 58880 45200
rect 1104 45126 2350 45178
rect 2402 45126 2414 45178
rect 2466 45126 2478 45178
rect 2530 45126 2542 45178
rect 2594 45126 2606 45178
rect 2658 45126 33070 45178
rect 33122 45126 33134 45178
rect 33186 45126 33198 45178
rect 33250 45126 33262 45178
rect 33314 45126 33326 45178
rect 33378 45126 58880 45178
rect 1104 45104 58880 45126
rect 58250 44888 58256 44940
rect 58308 44888 58314 44940
rect 58526 44820 58532 44872
rect 58584 44820 58590 44872
rect 1104 44634 58880 44656
rect 1104 44582 3010 44634
rect 3062 44582 3074 44634
rect 3126 44582 3138 44634
rect 3190 44582 3202 44634
rect 3254 44582 3266 44634
rect 3318 44582 33730 44634
rect 33782 44582 33794 44634
rect 33846 44582 33858 44634
rect 33910 44582 33922 44634
rect 33974 44582 33986 44634
rect 34038 44582 58880 44634
rect 1104 44560 58880 44582
rect 1104 44090 58880 44112
rect 1104 44038 2350 44090
rect 2402 44038 2414 44090
rect 2466 44038 2478 44090
rect 2530 44038 2542 44090
rect 2594 44038 2606 44090
rect 2658 44038 33070 44090
rect 33122 44038 33134 44090
rect 33186 44038 33198 44090
rect 33250 44038 33262 44090
rect 33314 44038 33326 44090
rect 33378 44038 58880 44090
rect 1104 44016 58880 44038
rect 1104 43546 58880 43568
rect 1104 43494 3010 43546
rect 3062 43494 3074 43546
rect 3126 43494 3138 43546
rect 3190 43494 3202 43546
rect 3254 43494 3266 43546
rect 3318 43494 33730 43546
rect 33782 43494 33794 43546
rect 33846 43494 33858 43546
rect 33910 43494 33922 43546
rect 33974 43494 33986 43546
rect 34038 43494 58880 43546
rect 1104 43472 58880 43494
rect 1104 43002 58880 43024
rect 1104 42950 2350 43002
rect 2402 42950 2414 43002
rect 2466 42950 2478 43002
rect 2530 42950 2542 43002
rect 2594 42950 2606 43002
rect 2658 42950 33070 43002
rect 33122 42950 33134 43002
rect 33186 42950 33198 43002
rect 33250 42950 33262 43002
rect 33314 42950 33326 43002
rect 33378 42950 58880 43002
rect 1104 42928 58880 42950
rect 1104 42458 58880 42480
rect 1104 42406 3010 42458
rect 3062 42406 3074 42458
rect 3126 42406 3138 42458
rect 3190 42406 3202 42458
rect 3254 42406 3266 42458
rect 3318 42406 33730 42458
rect 33782 42406 33794 42458
rect 33846 42406 33858 42458
rect 33910 42406 33922 42458
rect 33974 42406 33986 42458
rect 34038 42406 58880 42458
rect 1104 42384 58880 42406
rect 1104 41914 58880 41936
rect 1104 41862 2350 41914
rect 2402 41862 2414 41914
rect 2466 41862 2478 41914
rect 2530 41862 2542 41914
rect 2594 41862 2606 41914
rect 2658 41862 33070 41914
rect 33122 41862 33134 41914
rect 33186 41862 33198 41914
rect 33250 41862 33262 41914
rect 33314 41862 33326 41914
rect 33378 41862 58880 41914
rect 1104 41840 58880 41862
rect 1104 41370 58880 41392
rect 1104 41318 3010 41370
rect 3062 41318 3074 41370
rect 3126 41318 3138 41370
rect 3190 41318 3202 41370
rect 3254 41318 3266 41370
rect 3318 41318 33730 41370
rect 33782 41318 33794 41370
rect 33846 41318 33858 41370
rect 33910 41318 33922 41370
rect 33974 41318 33986 41370
rect 34038 41318 58880 41370
rect 1104 41296 58880 41318
rect 1104 40826 58880 40848
rect 1104 40774 2350 40826
rect 2402 40774 2414 40826
rect 2466 40774 2478 40826
rect 2530 40774 2542 40826
rect 2594 40774 2606 40826
rect 2658 40774 33070 40826
rect 33122 40774 33134 40826
rect 33186 40774 33198 40826
rect 33250 40774 33262 40826
rect 33314 40774 33326 40826
rect 33378 40774 58880 40826
rect 1104 40752 58880 40774
rect 1104 40282 58880 40304
rect 1104 40230 3010 40282
rect 3062 40230 3074 40282
rect 3126 40230 3138 40282
rect 3190 40230 3202 40282
rect 3254 40230 3266 40282
rect 3318 40230 33730 40282
rect 33782 40230 33794 40282
rect 33846 40230 33858 40282
rect 33910 40230 33922 40282
rect 33974 40230 33986 40282
rect 34038 40230 58880 40282
rect 1104 40208 58880 40230
rect 1104 39738 58880 39760
rect 1104 39686 2350 39738
rect 2402 39686 2414 39738
rect 2466 39686 2478 39738
rect 2530 39686 2542 39738
rect 2594 39686 2606 39738
rect 2658 39686 33070 39738
rect 33122 39686 33134 39738
rect 33186 39686 33198 39738
rect 33250 39686 33262 39738
rect 33314 39686 33326 39738
rect 33378 39686 58880 39738
rect 1104 39664 58880 39686
rect 1104 39194 58880 39216
rect 1104 39142 3010 39194
rect 3062 39142 3074 39194
rect 3126 39142 3138 39194
rect 3190 39142 3202 39194
rect 3254 39142 3266 39194
rect 3318 39142 33730 39194
rect 33782 39142 33794 39194
rect 33846 39142 33858 39194
rect 33910 39142 33922 39194
rect 33974 39142 33986 39194
rect 34038 39142 58880 39194
rect 1104 39120 58880 39142
rect 1104 38650 58880 38672
rect 1104 38598 2350 38650
rect 2402 38598 2414 38650
rect 2466 38598 2478 38650
rect 2530 38598 2542 38650
rect 2594 38598 2606 38650
rect 2658 38598 33070 38650
rect 33122 38598 33134 38650
rect 33186 38598 33198 38650
rect 33250 38598 33262 38650
rect 33314 38598 33326 38650
rect 33378 38598 58880 38650
rect 1104 38576 58880 38598
rect 1104 38106 58880 38128
rect 1104 38054 3010 38106
rect 3062 38054 3074 38106
rect 3126 38054 3138 38106
rect 3190 38054 3202 38106
rect 3254 38054 3266 38106
rect 3318 38054 33730 38106
rect 33782 38054 33794 38106
rect 33846 38054 33858 38106
rect 33910 38054 33922 38106
rect 33974 38054 33986 38106
rect 34038 38054 58880 38106
rect 1104 38032 58880 38054
rect 1104 37562 58880 37584
rect 1104 37510 2350 37562
rect 2402 37510 2414 37562
rect 2466 37510 2478 37562
rect 2530 37510 2542 37562
rect 2594 37510 2606 37562
rect 2658 37510 33070 37562
rect 33122 37510 33134 37562
rect 33186 37510 33198 37562
rect 33250 37510 33262 37562
rect 33314 37510 33326 37562
rect 33378 37510 58880 37562
rect 1104 37488 58880 37510
rect 1104 37018 58880 37040
rect 1104 36966 3010 37018
rect 3062 36966 3074 37018
rect 3126 36966 3138 37018
rect 3190 36966 3202 37018
rect 3254 36966 3266 37018
rect 3318 36966 33730 37018
rect 33782 36966 33794 37018
rect 33846 36966 33858 37018
rect 33910 36966 33922 37018
rect 33974 36966 33986 37018
rect 34038 36966 58880 37018
rect 1104 36944 58880 36966
rect 1104 36474 58880 36496
rect 1104 36422 2350 36474
rect 2402 36422 2414 36474
rect 2466 36422 2478 36474
rect 2530 36422 2542 36474
rect 2594 36422 2606 36474
rect 2658 36422 33070 36474
rect 33122 36422 33134 36474
rect 33186 36422 33198 36474
rect 33250 36422 33262 36474
rect 33314 36422 33326 36474
rect 33378 36422 58880 36474
rect 1104 36400 58880 36422
rect 1104 35930 58880 35952
rect 1104 35878 3010 35930
rect 3062 35878 3074 35930
rect 3126 35878 3138 35930
rect 3190 35878 3202 35930
rect 3254 35878 3266 35930
rect 3318 35878 33730 35930
rect 33782 35878 33794 35930
rect 33846 35878 33858 35930
rect 33910 35878 33922 35930
rect 33974 35878 33986 35930
rect 34038 35878 58880 35930
rect 1104 35856 58880 35878
rect 1104 35386 58880 35408
rect 1104 35334 2350 35386
rect 2402 35334 2414 35386
rect 2466 35334 2478 35386
rect 2530 35334 2542 35386
rect 2594 35334 2606 35386
rect 2658 35334 33070 35386
rect 33122 35334 33134 35386
rect 33186 35334 33198 35386
rect 33250 35334 33262 35386
rect 33314 35334 33326 35386
rect 33378 35334 58880 35386
rect 1104 35312 58880 35334
rect 1104 34842 58880 34864
rect 1104 34790 3010 34842
rect 3062 34790 3074 34842
rect 3126 34790 3138 34842
rect 3190 34790 3202 34842
rect 3254 34790 3266 34842
rect 3318 34790 33730 34842
rect 33782 34790 33794 34842
rect 33846 34790 33858 34842
rect 33910 34790 33922 34842
rect 33974 34790 33986 34842
rect 34038 34790 58880 34842
rect 1104 34768 58880 34790
rect 1104 34298 58880 34320
rect 1104 34246 2350 34298
rect 2402 34246 2414 34298
rect 2466 34246 2478 34298
rect 2530 34246 2542 34298
rect 2594 34246 2606 34298
rect 2658 34246 33070 34298
rect 33122 34246 33134 34298
rect 33186 34246 33198 34298
rect 33250 34246 33262 34298
rect 33314 34246 33326 34298
rect 33378 34246 58880 34298
rect 1104 34224 58880 34246
rect 1104 33754 58880 33776
rect 1104 33702 3010 33754
rect 3062 33702 3074 33754
rect 3126 33702 3138 33754
rect 3190 33702 3202 33754
rect 3254 33702 3266 33754
rect 3318 33702 33730 33754
rect 33782 33702 33794 33754
rect 33846 33702 33858 33754
rect 33910 33702 33922 33754
rect 33974 33702 33986 33754
rect 34038 33702 58880 33754
rect 1104 33680 58880 33702
rect 1104 33210 58880 33232
rect 1104 33158 2350 33210
rect 2402 33158 2414 33210
rect 2466 33158 2478 33210
rect 2530 33158 2542 33210
rect 2594 33158 2606 33210
rect 2658 33158 33070 33210
rect 33122 33158 33134 33210
rect 33186 33158 33198 33210
rect 33250 33158 33262 33210
rect 33314 33158 33326 33210
rect 33378 33158 58880 33210
rect 1104 33136 58880 33158
rect 1104 32666 58880 32688
rect 1104 32614 3010 32666
rect 3062 32614 3074 32666
rect 3126 32614 3138 32666
rect 3190 32614 3202 32666
rect 3254 32614 3266 32666
rect 3318 32614 33730 32666
rect 33782 32614 33794 32666
rect 33846 32614 33858 32666
rect 33910 32614 33922 32666
rect 33974 32614 33986 32666
rect 34038 32614 58880 32666
rect 1104 32592 58880 32614
rect 1104 32122 58880 32144
rect 1104 32070 2350 32122
rect 2402 32070 2414 32122
rect 2466 32070 2478 32122
rect 2530 32070 2542 32122
rect 2594 32070 2606 32122
rect 2658 32070 33070 32122
rect 33122 32070 33134 32122
rect 33186 32070 33198 32122
rect 33250 32070 33262 32122
rect 33314 32070 33326 32122
rect 33378 32070 58880 32122
rect 1104 32048 58880 32070
rect 1104 31578 58880 31600
rect 1104 31526 3010 31578
rect 3062 31526 3074 31578
rect 3126 31526 3138 31578
rect 3190 31526 3202 31578
rect 3254 31526 3266 31578
rect 3318 31526 33730 31578
rect 33782 31526 33794 31578
rect 33846 31526 33858 31578
rect 33910 31526 33922 31578
rect 33974 31526 33986 31578
rect 34038 31526 58880 31578
rect 1104 31504 58880 31526
rect 1104 31034 58880 31056
rect 1104 30982 2350 31034
rect 2402 30982 2414 31034
rect 2466 30982 2478 31034
rect 2530 30982 2542 31034
rect 2594 30982 2606 31034
rect 2658 30982 33070 31034
rect 33122 30982 33134 31034
rect 33186 30982 33198 31034
rect 33250 30982 33262 31034
rect 33314 30982 33326 31034
rect 33378 30982 58880 31034
rect 1104 30960 58880 30982
rect 1104 30490 58880 30512
rect 1104 30438 3010 30490
rect 3062 30438 3074 30490
rect 3126 30438 3138 30490
rect 3190 30438 3202 30490
rect 3254 30438 3266 30490
rect 3318 30438 33730 30490
rect 33782 30438 33794 30490
rect 33846 30438 33858 30490
rect 33910 30438 33922 30490
rect 33974 30438 33986 30490
rect 34038 30438 58880 30490
rect 1104 30416 58880 30438
rect 1104 29946 58880 29968
rect 1104 29894 2350 29946
rect 2402 29894 2414 29946
rect 2466 29894 2478 29946
rect 2530 29894 2542 29946
rect 2594 29894 2606 29946
rect 2658 29894 33070 29946
rect 33122 29894 33134 29946
rect 33186 29894 33198 29946
rect 33250 29894 33262 29946
rect 33314 29894 33326 29946
rect 33378 29894 58880 29946
rect 1104 29872 58880 29894
rect 1104 29402 58880 29424
rect 1104 29350 3010 29402
rect 3062 29350 3074 29402
rect 3126 29350 3138 29402
rect 3190 29350 3202 29402
rect 3254 29350 3266 29402
rect 3318 29350 33730 29402
rect 33782 29350 33794 29402
rect 33846 29350 33858 29402
rect 33910 29350 33922 29402
rect 33974 29350 33986 29402
rect 34038 29350 58880 29402
rect 1104 29328 58880 29350
rect 1104 28858 58880 28880
rect 1104 28806 2350 28858
rect 2402 28806 2414 28858
rect 2466 28806 2478 28858
rect 2530 28806 2542 28858
rect 2594 28806 2606 28858
rect 2658 28806 33070 28858
rect 33122 28806 33134 28858
rect 33186 28806 33198 28858
rect 33250 28806 33262 28858
rect 33314 28806 33326 28858
rect 33378 28806 58880 28858
rect 1104 28784 58880 28806
rect 1104 28314 58880 28336
rect 1104 28262 3010 28314
rect 3062 28262 3074 28314
rect 3126 28262 3138 28314
rect 3190 28262 3202 28314
rect 3254 28262 3266 28314
rect 3318 28262 33730 28314
rect 33782 28262 33794 28314
rect 33846 28262 33858 28314
rect 33910 28262 33922 28314
rect 33974 28262 33986 28314
rect 34038 28262 58880 28314
rect 1104 28240 58880 28262
rect 1104 27770 58880 27792
rect 1104 27718 2350 27770
rect 2402 27718 2414 27770
rect 2466 27718 2478 27770
rect 2530 27718 2542 27770
rect 2594 27718 2606 27770
rect 2658 27718 33070 27770
rect 33122 27718 33134 27770
rect 33186 27718 33198 27770
rect 33250 27718 33262 27770
rect 33314 27718 33326 27770
rect 33378 27718 58880 27770
rect 1104 27696 58880 27718
rect 1104 27226 58880 27248
rect 1104 27174 3010 27226
rect 3062 27174 3074 27226
rect 3126 27174 3138 27226
rect 3190 27174 3202 27226
rect 3254 27174 3266 27226
rect 3318 27174 33730 27226
rect 33782 27174 33794 27226
rect 33846 27174 33858 27226
rect 33910 27174 33922 27226
rect 33974 27174 33986 27226
rect 34038 27174 58880 27226
rect 1104 27152 58880 27174
rect 1104 26682 58880 26704
rect 1104 26630 2350 26682
rect 2402 26630 2414 26682
rect 2466 26630 2478 26682
rect 2530 26630 2542 26682
rect 2594 26630 2606 26682
rect 2658 26630 33070 26682
rect 33122 26630 33134 26682
rect 33186 26630 33198 26682
rect 33250 26630 33262 26682
rect 33314 26630 33326 26682
rect 33378 26630 58880 26682
rect 1104 26608 58880 26630
rect 1104 26138 58880 26160
rect 1104 26086 3010 26138
rect 3062 26086 3074 26138
rect 3126 26086 3138 26138
rect 3190 26086 3202 26138
rect 3254 26086 3266 26138
rect 3318 26086 33730 26138
rect 33782 26086 33794 26138
rect 33846 26086 33858 26138
rect 33910 26086 33922 26138
rect 33974 26086 33986 26138
rect 34038 26086 58880 26138
rect 1104 26064 58880 26086
rect 1104 25594 58880 25616
rect 1104 25542 2350 25594
rect 2402 25542 2414 25594
rect 2466 25542 2478 25594
rect 2530 25542 2542 25594
rect 2594 25542 2606 25594
rect 2658 25542 33070 25594
rect 33122 25542 33134 25594
rect 33186 25542 33198 25594
rect 33250 25542 33262 25594
rect 33314 25542 33326 25594
rect 33378 25542 58880 25594
rect 1104 25520 58880 25542
rect 1104 25050 58880 25072
rect 1104 24998 3010 25050
rect 3062 24998 3074 25050
rect 3126 24998 3138 25050
rect 3190 24998 3202 25050
rect 3254 24998 3266 25050
rect 3318 24998 33730 25050
rect 33782 24998 33794 25050
rect 33846 24998 33858 25050
rect 33910 24998 33922 25050
rect 33974 24998 33986 25050
rect 34038 24998 58880 25050
rect 1104 24976 58880 24998
rect 1104 24506 58880 24528
rect 1104 24454 2350 24506
rect 2402 24454 2414 24506
rect 2466 24454 2478 24506
rect 2530 24454 2542 24506
rect 2594 24454 2606 24506
rect 2658 24454 33070 24506
rect 33122 24454 33134 24506
rect 33186 24454 33198 24506
rect 33250 24454 33262 24506
rect 33314 24454 33326 24506
rect 33378 24454 58880 24506
rect 1104 24432 58880 24454
rect 1104 23962 58880 23984
rect 1104 23910 3010 23962
rect 3062 23910 3074 23962
rect 3126 23910 3138 23962
rect 3190 23910 3202 23962
rect 3254 23910 3266 23962
rect 3318 23910 33730 23962
rect 33782 23910 33794 23962
rect 33846 23910 33858 23962
rect 33910 23910 33922 23962
rect 33974 23910 33986 23962
rect 34038 23910 58880 23962
rect 1104 23888 58880 23910
rect 1104 23418 58880 23440
rect 1104 23366 2350 23418
rect 2402 23366 2414 23418
rect 2466 23366 2478 23418
rect 2530 23366 2542 23418
rect 2594 23366 2606 23418
rect 2658 23366 33070 23418
rect 33122 23366 33134 23418
rect 33186 23366 33198 23418
rect 33250 23366 33262 23418
rect 33314 23366 33326 23418
rect 33378 23366 58880 23418
rect 1104 23344 58880 23366
rect 1104 22874 58880 22896
rect 1104 22822 3010 22874
rect 3062 22822 3074 22874
rect 3126 22822 3138 22874
rect 3190 22822 3202 22874
rect 3254 22822 3266 22874
rect 3318 22822 33730 22874
rect 33782 22822 33794 22874
rect 33846 22822 33858 22874
rect 33910 22822 33922 22874
rect 33974 22822 33986 22874
rect 34038 22822 58880 22874
rect 1104 22800 58880 22822
rect 1104 22330 58880 22352
rect 1104 22278 2350 22330
rect 2402 22278 2414 22330
rect 2466 22278 2478 22330
rect 2530 22278 2542 22330
rect 2594 22278 2606 22330
rect 2658 22278 33070 22330
rect 33122 22278 33134 22330
rect 33186 22278 33198 22330
rect 33250 22278 33262 22330
rect 33314 22278 33326 22330
rect 33378 22278 58880 22330
rect 1104 22256 58880 22278
rect 1104 21786 58880 21808
rect 1104 21734 3010 21786
rect 3062 21734 3074 21786
rect 3126 21734 3138 21786
rect 3190 21734 3202 21786
rect 3254 21734 3266 21786
rect 3318 21734 33730 21786
rect 33782 21734 33794 21786
rect 33846 21734 33858 21786
rect 33910 21734 33922 21786
rect 33974 21734 33986 21786
rect 34038 21734 58880 21786
rect 1104 21712 58880 21734
rect 1104 21242 58880 21264
rect 1104 21190 2350 21242
rect 2402 21190 2414 21242
rect 2466 21190 2478 21242
rect 2530 21190 2542 21242
rect 2594 21190 2606 21242
rect 2658 21190 33070 21242
rect 33122 21190 33134 21242
rect 33186 21190 33198 21242
rect 33250 21190 33262 21242
rect 33314 21190 33326 21242
rect 33378 21190 58880 21242
rect 1104 21168 58880 21190
rect 1104 20698 58880 20720
rect 1104 20646 3010 20698
rect 3062 20646 3074 20698
rect 3126 20646 3138 20698
rect 3190 20646 3202 20698
rect 3254 20646 3266 20698
rect 3318 20646 33730 20698
rect 33782 20646 33794 20698
rect 33846 20646 33858 20698
rect 33910 20646 33922 20698
rect 33974 20646 33986 20698
rect 34038 20646 58880 20698
rect 1104 20624 58880 20646
rect 1104 20154 58880 20176
rect 1104 20102 2350 20154
rect 2402 20102 2414 20154
rect 2466 20102 2478 20154
rect 2530 20102 2542 20154
rect 2594 20102 2606 20154
rect 2658 20102 33070 20154
rect 33122 20102 33134 20154
rect 33186 20102 33198 20154
rect 33250 20102 33262 20154
rect 33314 20102 33326 20154
rect 33378 20102 58880 20154
rect 1104 20080 58880 20102
rect 1104 19610 58880 19632
rect 1104 19558 3010 19610
rect 3062 19558 3074 19610
rect 3126 19558 3138 19610
rect 3190 19558 3202 19610
rect 3254 19558 3266 19610
rect 3318 19558 33730 19610
rect 33782 19558 33794 19610
rect 33846 19558 33858 19610
rect 33910 19558 33922 19610
rect 33974 19558 33986 19610
rect 34038 19558 58880 19610
rect 1104 19536 58880 19558
rect 1104 19066 58880 19088
rect 1104 19014 2350 19066
rect 2402 19014 2414 19066
rect 2466 19014 2478 19066
rect 2530 19014 2542 19066
rect 2594 19014 2606 19066
rect 2658 19014 33070 19066
rect 33122 19014 33134 19066
rect 33186 19014 33198 19066
rect 33250 19014 33262 19066
rect 33314 19014 33326 19066
rect 33378 19014 58880 19066
rect 1104 18992 58880 19014
rect 1104 18522 58880 18544
rect 1104 18470 3010 18522
rect 3062 18470 3074 18522
rect 3126 18470 3138 18522
rect 3190 18470 3202 18522
rect 3254 18470 3266 18522
rect 3318 18470 33730 18522
rect 33782 18470 33794 18522
rect 33846 18470 33858 18522
rect 33910 18470 33922 18522
rect 33974 18470 33986 18522
rect 34038 18470 58880 18522
rect 1104 18448 58880 18470
rect 1104 17978 58880 18000
rect 1104 17926 2350 17978
rect 2402 17926 2414 17978
rect 2466 17926 2478 17978
rect 2530 17926 2542 17978
rect 2594 17926 2606 17978
rect 2658 17926 33070 17978
rect 33122 17926 33134 17978
rect 33186 17926 33198 17978
rect 33250 17926 33262 17978
rect 33314 17926 33326 17978
rect 33378 17926 58880 17978
rect 1104 17904 58880 17926
rect 1104 17434 58880 17456
rect 1104 17382 3010 17434
rect 3062 17382 3074 17434
rect 3126 17382 3138 17434
rect 3190 17382 3202 17434
rect 3254 17382 3266 17434
rect 3318 17382 33730 17434
rect 33782 17382 33794 17434
rect 33846 17382 33858 17434
rect 33910 17382 33922 17434
rect 33974 17382 33986 17434
rect 34038 17382 58880 17434
rect 1104 17360 58880 17382
rect 1104 16890 58880 16912
rect 1104 16838 2350 16890
rect 2402 16838 2414 16890
rect 2466 16838 2478 16890
rect 2530 16838 2542 16890
rect 2594 16838 2606 16890
rect 2658 16838 33070 16890
rect 33122 16838 33134 16890
rect 33186 16838 33198 16890
rect 33250 16838 33262 16890
rect 33314 16838 33326 16890
rect 33378 16838 58880 16890
rect 1104 16816 58880 16838
rect 1104 16346 58880 16368
rect 1104 16294 3010 16346
rect 3062 16294 3074 16346
rect 3126 16294 3138 16346
rect 3190 16294 3202 16346
rect 3254 16294 3266 16346
rect 3318 16294 33730 16346
rect 33782 16294 33794 16346
rect 33846 16294 33858 16346
rect 33910 16294 33922 16346
rect 33974 16294 33986 16346
rect 34038 16294 58880 16346
rect 1104 16272 58880 16294
rect 1104 15802 58880 15824
rect 1104 15750 2350 15802
rect 2402 15750 2414 15802
rect 2466 15750 2478 15802
rect 2530 15750 2542 15802
rect 2594 15750 2606 15802
rect 2658 15750 33070 15802
rect 33122 15750 33134 15802
rect 33186 15750 33198 15802
rect 33250 15750 33262 15802
rect 33314 15750 33326 15802
rect 33378 15750 58880 15802
rect 1104 15728 58880 15750
rect 1104 15258 58880 15280
rect 1104 15206 3010 15258
rect 3062 15206 3074 15258
rect 3126 15206 3138 15258
rect 3190 15206 3202 15258
rect 3254 15206 3266 15258
rect 3318 15206 33730 15258
rect 33782 15206 33794 15258
rect 33846 15206 33858 15258
rect 33910 15206 33922 15258
rect 33974 15206 33986 15258
rect 34038 15206 58880 15258
rect 1104 15184 58880 15206
rect 38010 15104 38016 15156
rect 38068 15144 38074 15156
rect 56502 15144 56508 15156
rect 38068 15116 56508 15144
rect 38068 15104 38074 15116
rect 56502 15104 56508 15116
rect 56560 15104 56566 15156
rect 1104 14714 58880 14736
rect 1104 14662 2350 14714
rect 2402 14662 2414 14714
rect 2466 14662 2478 14714
rect 2530 14662 2542 14714
rect 2594 14662 2606 14714
rect 2658 14662 33070 14714
rect 33122 14662 33134 14714
rect 33186 14662 33198 14714
rect 33250 14662 33262 14714
rect 33314 14662 33326 14714
rect 33378 14662 58880 14714
rect 1104 14640 58880 14662
rect 1104 14170 58880 14192
rect 1104 14118 3010 14170
rect 3062 14118 3074 14170
rect 3126 14118 3138 14170
rect 3190 14118 3202 14170
rect 3254 14118 3266 14170
rect 3318 14118 33730 14170
rect 33782 14118 33794 14170
rect 33846 14118 33858 14170
rect 33910 14118 33922 14170
rect 33974 14118 33986 14170
rect 34038 14118 58880 14170
rect 1104 14096 58880 14118
rect 1104 13626 58880 13648
rect 1104 13574 2350 13626
rect 2402 13574 2414 13626
rect 2466 13574 2478 13626
rect 2530 13574 2542 13626
rect 2594 13574 2606 13626
rect 2658 13574 33070 13626
rect 33122 13574 33134 13626
rect 33186 13574 33198 13626
rect 33250 13574 33262 13626
rect 33314 13574 33326 13626
rect 33378 13574 58880 13626
rect 1104 13552 58880 13574
rect 1104 13082 58880 13104
rect 1104 13030 3010 13082
rect 3062 13030 3074 13082
rect 3126 13030 3138 13082
rect 3190 13030 3202 13082
rect 3254 13030 3266 13082
rect 3318 13030 33730 13082
rect 33782 13030 33794 13082
rect 33846 13030 33858 13082
rect 33910 13030 33922 13082
rect 33974 13030 33986 13082
rect 34038 13030 58880 13082
rect 1104 13008 58880 13030
rect 1104 12538 58880 12560
rect 1104 12486 2350 12538
rect 2402 12486 2414 12538
rect 2466 12486 2478 12538
rect 2530 12486 2542 12538
rect 2594 12486 2606 12538
rect 2658 12486 33070 12538
rect 33122 12486 33134 12538
rect 33186 12486 33198 12538
rect 33250 12486 33262 12538
rect 33314 12486 33326 12538
rect 33378 12486 58880 12538
rect 1104 12464 58880 12486
rect 1104 11994 58880 12016
rect 1104 11942 3010 11994
rect 3062 11942 3074 11994
rect 3126 11942 3138 11994
rect 3190 11942 3202 11994
rect 3254 11942 3266 11994
rect 3318 11942 33730 11994
rect 33782 11942 33794 11994
rect 33846 11942 33858 11994
rect 33910 11942 33922 11994
rect 33974 11942 33986 11994
rect 34038 11942 58880 11994
rect 1104 11920 58880 11942
rect 1104 11450 58880 11472
rect 1104 11398 2350 11450
rect 2402 11398 2414 11450
rect 2466 11398 2478 11450
rect 2530 11398 2542 11450
rect 2594 11398 2606 11450
rect 2658 11398 33070 11450
rect 33122 11398 33134 11450
rect 33186 11398 33198 11450
rect 33250 11398 33262 11450
rect 33314 11398 33326 11450
rect 33378 11398 58880 11450
rect 1104 11376 58880 11398
rect 1104 10906 58880 10928
rect 1104 10854 3010 10906
rect 3062 10854 3074 10906
rect 3126 10854 3138 10906
rect 3190 10854 3202 10906
rect 3254 10854 3266 10906
rect 3318 10854 33730 10906
rect 33782 10854 33794 10906
rect 33846 10854 33858 10906
rect 33910 10854 33922 10906
rect 33974 10854 33986 10906
rect 34038 10854 58880 10906
rect 1104 10832 58880 10854
rect 1104 10362 58880 10384
rect 1104 10310 2350 10362
rect 2402 10310 2414 10362
rect 2466 10310 2478 10362
rect 2530 10310 2542 10362
rect 2594 10310 2606 10362
rect 2658 10310 33070 10362
rect 33122 10310 33134 10362
rect 33186 10310 33198 10362
rect 33250 10310 33262 10362
rect 33314 10310 33326 10362
rect 33378 10310 58880 10362
rect 1104 10288 58880 10310
rect 1104 9818 58880 9840
rect 1104 9766 3010 9818
rect 3062 9766 3074 9818
rect 3126 9766 3138 9818
rect 3190 9766 3202 9818
rect 3254 9766 3266 9818
rect 3318 9766 33730 9818
rect 33782 9766 33794 9818
rect 33846 9766 33858 9818
rect 33910 9766 33922 9818
rect 33974 9766 33986 9818
rect 34038 9766 58880 9818
rect 1104 9744 58880 9766
rect 1104 9274 58880 9296
rect 1104 9222 2350 9274
rect 2402 9222 2414 9274
rect 2466 9222 2478 9274
rect 2530 9222 2542 9274
rect 2594 9222 2606 9274
rect 2658 9222 33070 9274
rect 33122 9222 33134 9274
rect 33186 9222 33198 9274
rect 33250 9222 33262 9274
rect 33314 9222 33326 9274
rect 33378 9222 58880 9274
rect 1104 9200 58880 9222
rect 1104 8730 58880 8752
rect 1104 8678 3010 8730
rect 3062 8678 3074 8730
rect 3126 8678 3138 8730
rect 3190 8678 3202 8730
rect 3254 8678 3266 8730
rect 3318 8678 33730 8730
rect 33782 8678 33794 8730
rect 33846 8678 33858 8730
rect 33910 8678 33922 8730
rect 33974 8678 33986 8730
rect 34038 8678 58880 8730
rect 1104 8656 58880 8678
rect 1104 8186 58880 8208
rect 1104 8134 2350 8186
rect 2402 8134 2414 8186
rect 2466 8134 2478 8186
rect 2530 8134 2542 8186
rect 2594 8134 2606 8186
rect 2658 8134 33070 8186
rect 33122 8134 33134 8186
rect 33186 8134 33198 8186
rect 33250 8134 33262 8186
rect 33314 8134 33326 8186
rect 33378 8134 58880 8186
rect 1104 8112 58880 8134
rect 1104 7642 58880 7664
rect 1104 7590 3010 7642
rect 3062 7590 3074 7642
rect 3126 7590 3138 7642
rect 3190 7590 3202 7642
rect 3254 7590 3266 7642
rect 3318 7590 33730 7642
rect 33782 7590 33794 7642
rect 33846 7590 33858 7642
rect 33910 7590 33922 7642
rect 33974 7590 33986 7642
rect 34038 7590 58880 7642
rect 1104 7568 58880 7590
rect 1104 7098 58880 7120
rect 1104 7046 2350 7098
rect 2402 7046 2414 7098
rect 2466 7046 2478 7098
rect 2530 7046 2542 7098
rect 2594 7046 2606 7098
rect 2658 7046 33070 7098
rect 33122 7046 33134 7098
rect 33186 7046 33198 7098
rect 33250 7046 33262 7098
rect 33314 7046 33326 7098
rect 33378 7046 58880 7098
rect 1104 7024 58880 7046
rect 1104 6554 58880 6576
rect 1104 6502 3010 6554
rect 3062 6502 3074 6554
rect 3126 6502 3138 6554
rect 3190 6502 3202 6554
rect 3254 6502 3266 6554
rect 3318 6502 33730 6554
rect 33782 6502 33794 6554
rect 33846 6502 33858 6554
rect 33910 6502 33922 6554
rect 33974 6502 33986 6554
rect 34038 6502 58880 6554
rect 1104 6480 58880 6502
rect 1104 6010 58880 6032
rect 1104 5958 2350 6010
rect 2402 5958 2414 6010
rect 2466 5958 2478 6010
rect 2530 5958 2542 6010
rect 2594 5958 2606 6010
rect 2658 5958 33070 6010
rect 33122 5958 33134 6010
rect 33186 5958 33198 6010
rect 33250 5958 33262 6010
rect 33314 5958 33326 6010
rect 33378 5958 58880 6010
rect 1104 5936 58880 5958
rect 1104 5466 58880 5488
rect 1104 5414 3010 5466
rect 3062 5414 3074 5466
rect 3126 5414 3138 5466
rect 3190 5414 3202 5466
rect 3254 5414 3266 5466
rect 3318 5414 33730 5466
rect 33782 5414 33794 5466
rect 33846 5414 33858 5466
rect 33910 5414 33922 5466
rect 33974 5414 33986 5466
rect 34038 5414 58880 5466
rect 1104 5392 58880 5414
rect 1104 4922 58880 4944
rect 1104 4870 2350 4922
rect 2402 4870 2414 4922
rect 2466 4870 2478 4922
rect 2530 4870 2542 4922
rect 2594 4870 2606 4922
rect 2658 4870 33070 4922
rect 33122 4870 33134 4922
rect 33186 4870 33198 4922
rect 33250 4870 33262 4922
rect 33314 4870 33326 4922
rect 33378 4870 58880 4922
rect 1104 4848 58880 4870
rect 1104 4378 58880 4400
rect 1104 4326 3010 4378
rect 3062 4326 3074 4378
rect 3126 4326 3138 4378
rect 3190 4326 3202 4378
rect 3254 4326 3266 4378
rect 3318 4326 33730 4378
rect 33782 4326 33794 4378
rect 33846 4326 33858 4378
rect 33910 4326 33922 4378
rect 33974 4326 33986 4378
rect 34038 4326 58880 4378
rect 1104 4304 58880 4326
rect 1104 3834 58880 3856
rect 1104 3782 2350 3834
rect 2402 3782 2414 3834
rect 2466 3782 2478 3834
rect 2530 3782 2542 3834
rect 2594 3782 2606 3834
rect 2658 3782 33070 3834
rect 33122 3782 33134 3834
rect 33186 3782 33198 3834
rect 33250 3782 33262 3834
rect 33314 3782 33326 3834
rect 33378 3782 58880 3834
rect 1104 3760 58880 3782
rect 1104 3290 58880 3312
rect 1104 3238 3010 3290
rect 3062 3238 3074 3290
rect 3126 3238 3138 3290
rect 3190 3238 3202 3290
rect 3254 3238 3266 3290
rect 3318 3238 33730 3290
rect 33782 3238 33794 3290
rect 33846 3238 33858 3290
rect 33910 3238 33922 3290
rect 33974 3238 33986 3290
rect 34038 3238 58880 3290
rect 1104 3216 58880 3238
rect 1104 2746 58880 2768
rect 1104 2694 2350 2746
rect 2402 2694 2414 2746
rect 2466 2694 2478 2746
rect 2530 2694 2542 2746
rect 2594 2694 2606 2746
rect 2658 2694 33070 2746
rect 33122 2694 33134 2746
rect 33186 2694 33198 2746
rect 33250 2694 33262 2746
rect 33314 2694 33326 2746
rect 33378 2694 58880 2746
rect 1104 2672 58880 2694
rect 1104 2202 58880 2224
rect 1104 2150 3010 2202
rect 3062 2150 3074 2202
rect 3126 2150 3138 2202
rect 3190 2150 3202 2202
rect 3254 2150 3266 2202
rect 3318 2150 33730 2202
rect 33782 2150 33794 2202
rect 33846 2150 33858 2202
rect 33910 2150 33922 2202
rect 33974 2150 33986 2202
rect 34038 2150 58880 2202
rect 1104 2128 58880 2150
<< via1 >>
rect 3010 57638 3062 57690
rect 3074 57638 3126 57690
rect 3138 57638 3190 57690
rect 3202 57638 3254 57690
rect 3266 57638 3318 57690
rect 33730 57638 33782 57690
rect 33794 57638 33846 57690
rect 33858 57638 33910 57690
rect 33922 57638 33974 57690
rect 33986 57638 34038 57690
rect 6736 57536 6788 57588
rect 2872 57468 2924 57520
rect 4804 57468 4856 57520
rect 8668 57468 8720 57520
rect 10600 57468 10652 57520
rect 15292 57536 15344 57588
rect 26240 57579 26292 57588
rect 26240 57545 26249 57579
rect 26249 57545 26283 57579
rect 26283 57545 26292 57579
rect 26240 57536 26292 57545
rect 27988 57536 28040 57588
rect 30380 57579 30432 57588
rect 30380 57545 30389 57579
rect 30389 57545 30423 57579
rect 30423 57545 30432 57579
rect 30380 57536 30432 57545
rect 34152 57579 34204 57588
rect 34152 57545 34161 57579
rect 34161 57545 34195 57579
rect 34195 57545 34204 57579
rect 34152 57536 34204 57545
rect 35716 57536 35768 57588
rect 45376 57536 45428 57588
rect 47308 57536 47360 57588
rect 49700 57579 49752 57588
rect 49700 57545 49709 57579
rect 49709 57545 49743 57579
rect 49743 57545 49752 57579
rect 49700 57536 49752 57545
rect 51172 57536 51224 57588
rect 53104 57536 53156 57588
rect 55036 57536 55088 57588
rect 56968 57536 57020 57588
rect 12532 57468 12584 57520
rect 940 57400 992 57452
rect 4068 57400 4120 57452
rect 5264 57443 5316 57452
rect 5264 57409 5273 57443
rect 5273 57409 5307 57443
rect 5307 57409 5316 57443
rect 5264 57400 5316 57409
rect 7196 57443 7248 57452
rect 7196 57409 7205 57443
rect 7205 57409 7239 57443
rect 7239 57409 7248 57443
rect 7196 57400 7248 57409
rect 14464 57468 14516 57520
rect 15200 57468 15252 57520
rect 16396 57468 16448 57520
rect 18328 57468 18380 57520
rect 20260 57468 20312 57520
rect 22192 57468 22244 57520
rect 24124 57468 24176 57520
rect 31852 57468 31904 57520
rect 37648 57468 37700 57520
rect 39580 57468 39632 57520
rect 41512 57468 41564 57520
rect 43444 57468 43496 57520
rect 53012 57468 53064 57520
rect 56140 57468 56192 57520
rect 58900 57468 58952 57520
rect 16764 57400 16816 57452
rect 17224 57400 17276 57452
rect 18880 57400 18932 57452
rect 20720 57443 20772 57452
rect 20720 57409 20729 57443
rect 20729 57409 20763 57443
rect 20763 57409 20772 57443
rect 20720 57400 20772 57409
rect 22468 57400 22520 57452
rect 24768 57443 24820 57452
rect 24768 57409 24777 57443
rect 24777 57409 24811 57443
rect 24811 57409 24820 57443
rect 24768 57400 24820 57409
rect 27068 57400 27120 57452
rect 27712 57400 27764 57452
rect 30104 57443 30156 57452
rect 30104 57409 30113 57443
rect 30113 57409 30147 57443
rect 30147 57409 30156 57443
rect 30104 57400 30156 57409
rect 32496 57443 32548 57452
rect 32496 57409 32505 57443
rect 32505 57409 32539 57443
rect 32539 57409 32548 57443
rect 32496 57400 32548 57409
rect 34244 57443 34296 57452
rect 34244 57409 34253 57443
rect 34253 57409 34287 57443
rect 34287 57409 34296 57443
rect 34244 57400 34296 57409
rect 35900 57400 35952 57452
rect 38108 57443 38160 57452
rect 38108 57409 38117 57443
rect 38117 57409 38151 57443
rect 38151 57409 38160 57443
rect 38108 57400 38160 57409
rect 40224 57443 40276 57452
rect 40224 57409 40233 57443
rect 40233 57409 40267 57443
rect 40267 57409 40276 57443
rect 40224 57400 40276 57409
rect 41972 57443 42024 57452
rect 41972 57409 41981 57443
rect 41981 57409 42015 57443
rect 42015 57409 42024 57443
rect 41972 57400 42024 57409
rect 43904 57443 43956 57452
rect 43904 57409 43913 57443
rect 43913 57409 43947 57443
rect 43947 57409 43956 57443
rect 43904 57400 43956 57409
rect 45560 57443 45612 57452
rect 45560 57409 45569 57443
rect 45569 57409 45603 57443
rect 45603 57409 45612 57443
rect 45560 57400 45612 57409
rect 47676 57443 47728 57452
rect 47676 57409 47685 57443
rect 47685 57409 47719 57443
rect 47719 57409 47728 57443
rect 47676 57400 47728 57409
rect 49424 57443 49476 57452
rect 49424 57409 49433 57443
rect 49433 57409 49467 57443
rect 49467 57409 49476 57443
rect 49424 57400 49476 57409
rect 51172 57400 51224 57452
rect 52000 57400 52052 57452
rect 55864 57400 55916 57452
rect 16120 57264 16172 57316
rect 16856 57332 16908 57384
rect 2350 57094 2402 57146
rect 2414 57094 2466 57146
rect 2478 57094 2530 57146
rect 2542 57094 2594 57146
rect 2606 57094 2658 57146
rect 33070 57094 33122 57146
rect 33134 57094 33186 57146
rect 33198 57094 33250 57146
rect 33262 57094 33314 57146
rect 33326 57094 33378 57146
rect 5264 56924 5316 56976
rect 16028 56992 16080 57044
rect 21272 56992 21324 57044
rect 51540 56992 51592 57044
rect 52276 56992 52328 57044
rect 16396 56899 16448 56908
rect 16396 56865 16405 56899
rect 16405 56865 16439 56899
rect 16439 56865 16448 56899
rect 16396 56856 16448 56865
rect 20812 56924 20864 56976
rect 51080 56924 51132 56976
rect 17132 56856 17184 56908
rect 17316 56856 17368 56908
rect 17868 56856 17920 56908
rect 51540 56856 51592 56908
rect 52000 56899 52052 56908
rect 52000 56865 52009 56899
rect 52009 56865 52043 56899
rect 52043 56865 52052 56899
rect 52000 56856 52052 56865
rect 53012 56899 53064 56908
rect 53012 56865 53021 56899
rect 53021 56865 53055 56899
rect 53055 56865 53064 56899
rect 53012 56856 53064 56865
rect 15936 56788 15988 56840
rect 16212 56831 16264 56840
rect 16212 56797 16221 56831
rect 16221 56797 16255 56831
rect 16255 56797 16264 56831
rect 16212 56788 16264 56797
rect 16672 56831 16724 56840
rect 16672 56797 16681 56831
rect 16681 56797 16715 56831
rect 16715 56797 16724 56831
rect 16672 56788 16724 56797
rect 16856 56788 16908 56840
rect 18144 56788 18196 56840
rect 7196 56720 7248 56772
rect 17960 56720 18012 56772
rect 19524 56788 19576 56840
rect 22192 56831 22244 56840
rect 22192 56797 22201 56831
rect 22201 56797 22235 56831
rect 22235 56797 22244 56831
rect 22192 56788 22244 56797
rect 22468 56788 22520 56840
rect 27068 56831 27120 56840
rect 27068 56797 27077 56831
rect 27077 56797 27111 56831
rect 27111 56797 27120 56831
rect 27068 56788 27120 56797
rect 27804 56831 27856 56840
rect 27804 56797 27813 56831
rect 27813 56797 27847 56831
rect 27847 56797 27856 56831
rect 27804 56788 27856 56797
rect 28172 56831 28224 56840
rect 28172 56797 28181 56831
rect 28181 56797 28215 56831
rect 28215 56797 28224 56831
rect 28172 56788 28224 56797
rect 52736 56788 52788 56840
rect 16028 56652 16080 56704
rect 16948 56695 17000 56704
rect 16948 56661 16957 56695
rect 16957 56661 16991 56695
rect 16991 56661 17000 56695
rect 16948 56652 17000 56661
rect 17132 56652 17184 56704
rect 17408 56695 17460 56704
rect 17408 56661 17417 56695
rect 17417 56661 17451 56695
rect 17451 56661 17460 56695
rect 17408 56652 17460 56661
rect 18604 56652 18656 56704
rect 20904 56720 20956 56772
rect 22560 56652 22612 56704
rect 23664 56695 23716 56704
rect 23664 56661 23673 56695
rect 23673 56661 23707 56695
rect 23707 56661 23716 56695
rect 23664 56652 23716 56661
rect 26516 56695 26568 56704
rect 26516 56661 26525 56695
rect 26525 56661 26559 56695
rect 26559 56661 26568 56695
rect 26516 56652 26568 56661
rect 27160 56652 27212 56704
rect 27896 56652 27948 56704
rect 51632 56695 51684 56704
rect 51632 56661 51641 56695
rect 51641 56661 51675 56695
rect 51675 56661 51684 56695
rect 51632 56652 51684 56661
rect 52460 56695 52512 56704
rect 52460 56661 52469 56695
rect 52469 56661 52503 56695
rect 52503 56661 52512 56695
rect 52460 56652 52512 56661
rect 52920 56695 52972 56704
rect 52920 56661 52929 56695
rect 52929 56661 52963 56695
rect 52963 56661 52972 56695
rect 52920 56652 52972 56661
rect 3010 56550 3062 56602
rect 3074 56550 3126 56602
rect 3138 56550 3190 56602
rect 3202 56550 3254 56602
rect 3266 56550 3318 56602
rect 33730 56550 33782 56602
rect 33794 56550 33846 56602
rect 33858 56550 33910 56602
rect 33922 56550 33974 56602
rect 33986 56550 34038 56602
rect 15200 56491 15252 56500
rect 15200 56457 15209 56491
rect 15209 56457 15243 56491
rect 15243 56457 15252 56491
rect 15200 56448 15252 56457
rect 15292 56491 15344 56500
rect 15292 56457 15301 56491
rect 15301 56457 15335 56491
rect 15335 56457 15344 56491
rect 15292 56448 15344 56457
rect 15936 56380 15988 56432
rect 16120 56423 16172 56432
rect 16120 56389 16129 56423
rect 16129 56389 16163 56423
rect 16163 56389 16172 56423
rect 16120 56380 16172 56389
rect 16764 56448 16816 56500
rect 17776 56448 17828 56500
rect 16856 56380 16908 56432
rect 19248 56448 19300 56500
rect 17224 56312 17276 56364
rect 16396 56244 16448 56296
rect 17316 56244 17368 56296
rect 18880 56312 18932 56364
rect 18696 56287 18748 56296
rect 17592 56176 17644 56228
rect 18696 56253 18705 56287
rect 18705 56253 18739 56287
rect 18739 56253 18748 56287
rect 18696 56244 18748 56253
rect 20904 56380 20956 56432
rect 21272 56380 21324 56432
rect 23664 56448 23716 56500
rect 19432 56355 19484 56364
rect 19432 56321 19441 56355
rect 19441 56321 19475 56355
rect 19475 56321 19484 56355
rect 19432 56312 19484 56321
rect 18880 56176 18932 56228
rect 19984 56244 20036 56296
rect 22468 56312 22520 56364
rect 19432 56176 19484 56228
rect 22284 56244 22336 56296
rect 23756 56380 23808 56432
rect 24768 56448 24820 56500
rect 26516 56448 26568 56500
rect 27804 56448 27856 56500
rect 28172 56491 28224 56500
rect 28172 56457 28181 56491
rect 28181 56457 28215 56491
rect 28215 56457 28224 56491
rect 28172 56448 28224 56457
rect 15660 56151 15712 56160
rect 15660 56117 15669 56151
rect 15669 56117 15703 56151
rect 15703 56117 15712 56151
rect 15660 56108 15712 56117
rect 16028 56108 16080 56160
rect 17500 56108 17552 56160
rect 18328 56108 18380 56160
rect 19340 56108 19392 56160
rect 19616 56108 19668 56160
rect 19708 56108 19760 56160
rect 19892 56151 19944 56160
rect 19892 56117 19901 56151
rect 19901 56117 19935 56151
rect 19935 56117 19944 56151
rect 19892 56108 19944 56117
rect 27068 56380 27120 56432
rect 27712 56423 27764 56432
rect 27160 56355 27212 56364
rect 27160 56321 27169 56355
rect 27169 56321 27203 56355
rect 27203 56321 27212 56355
rect 27160 56312 27212 56321
rect 27712 56389 27721 56423
rect 27721 56389 27755 56423
rect 27755 56389 27764 56423
rect 27712 56380 27764 56389
rect 30104 56380 30156 56432
rect 28724 56287 28776 56296
rect 28724 56253 28733 56287
rect 28733 56253 28767 56287
rect 28767 56253 28776 56287
rect 28724 56244 28776 56253
rect 32220 56448 32272 56500
rect 32496 56448 32548 56500
rect 35900 56448 35952 56500
rect 32220 56244 32272 56296
rect 32680 56287 32732 56296
rect 32680 56253 32689 56287
rect 32689 56253 32723 56287
rect 32723 56253 32732 56287
rect 32680 56244 32732 56253
rect 34244 56287 34296 56296
rect 34244 56253 34253 56287
rect 34253 56253 34287 56287
rect 34287 56253 34296 56287
rect 34244 56244 34296 56253
rect 36268 56312 36320 56364
rect 38108 56448 38160 56500
rect 40224 56448 40276 56500
rect 43904 56380 43956 56432
rect 46940 56380 46992 56432
rect 47676 56380 47728 56432
rect 41604 56244 41656 56296
rect 41972 56244 42024 56296
rect 43720 56287 43772 56296
rect 43720 56253 43729 56287
rect 43729 56253 43763 56287
rect 43763 56253 43772 56287
rect 43720 56244 43772 56253
rect 45836 56312 45888 56364
rect 49424 56448 49476 56500
rect 49792 56491 49844 56500
rect 49792 56457 49801 56491
rect 49801 56457 49835 56491
rect 49835 56457 49844 56491
rect 49792 56448 49844 56457
rect 52000 56448 52052 56500
rect 52552 56448 52604 56500
rect 52736 56491 52788 56500
rect 52736 56457 52745 56491
rect 52745 56457 52779 56491
rect 52779 56457 52788 56491
rect 52736 56448 52788 56457
rect 51172 56380 51224 56432
rect 52920 56380 52972 56432
rect 55220 56380 55272 56432
rect 55864 56380 55916 56432
rect 45008 56244 45060 56296
rect 49056 56287 49108 56296
rect 49056 56253 49065 56287
rect 49065 56253 49099 56287
rect 49099 56253 49108 56287
rect 49056 56244 49108 56253
rect 51080 56312 51132 56364
rect 20720 56108 20772 56160
rect 21824 56108 21876 56160
rect 22100 56108 22152 56160
rect 22376 56108 22428 56160
rect 22744 56108 22796 56160
rect 25044 56108 25096 56160
rect 26976 56151 27028 56160
rect 26976 56117 26985 56151
rect 26985 56117 27019 56151
rect 27019 56117 27028 56151
rect 26976 56108 27028 56117
rect 28080 56108 28132 56160
rect 32404 56108 32456 56160
rect 34796 56151 34848 56160
rect 34796 56117 34805 56151
rect 34805 56117 34839 56151
rect 34839 56117 34848 56151
rect 34796 56108 34848 56117
rect 37740 56108 37792 56160
rect 38660 56108 38712 56160
rect 40132 56108 40184 56160
rect 41972 56108 42024 56160
rect 43444 56108 43496 56160
rect 44364 56108 44416 56160
rect 44916 56151 44968 56160
rect 44916 56117 44925 56151
rect 44925 56117 44959 56151
rect 44959 56117 44968 56151
rect 44916 56108 44968 56117
rect 49056 56108 49108 56160
rect 51540 56244 51592 56296
rect 51724 56176 51776 56228
rect 52460 56312 52512 56364
rect 55312 56312 55364 56364
rect 56140 56312 56192 56364
rect 52276 56244 52328 56296
rect 51080 56108 51132 56160
rect 52000 56108 52052 56160
rect 2350 56006 2402 56058
rect 2414 56006 2466 56058
rect 2478 56006 2530 56058
rect 2542 56006 2594 56058
rect 2606 56006 2658 56058
rect 33070 56006 33122 56058
rect 33134 56006 33186 56058
rect 33198 56006 33250 56058
rect 33262 56006 33314 56058
rect 33326 56006 33378 56058
rect 16672 55904 16724 55956
rect 18144 55947 18196 55956
rect 18144 55913 18153 55947
rect 18153 55913 18187 55947
rect 18187 55913 18196 55947
rect 18144 55904 18196 55913
rect 18696 55904 18748 55956
rect 19800 55904 19852 55956
rect 22376 55904 22428 55956
rect 17868 55836 17920 55888
rect 19340 55836 19392 55888
rect 19616 55836 19668 55888
rect 20444 55836 20496 55888
rect 21916 55836 21968 55888
rect 23756 55836 23808 55888
rect 24676 55836 24728 55888
rect 27712 55836 27764 55888
rect 28724 55836 28776 55888
rect 43720 55904 43772 55956
rect 45008 55947 45060 55956
rect 45008 55913 45017 55947
rect 45017 55913 45051 55947
rect 45051 55913 45060 55947
rect 45008 55904 45060 55913
rect 32680 55836 32732 55888
rect 4068 55768 4120 55820
rect 15660 55700 15712 55752
rect 16028 55743 16080 55752
rect 16028 55709 16037 55743
rect 16037 55709 16071 55743
rect 16071 55709 16080 55743
rect 16028 55700 16080 55709
rect 16948 55700 17000 55752
rect 17316 55768 17368 55820
rect 17592 55811 17644 55820
rect 17592 55777 17601 55811
rect 17601 55777 17635 55811
rect 17635 55777 17644 55811
rect 17592 55768 17644 55777
rect 17224 55700 17276 55752
rect 16120 55632 16172 55684
rect 18604 55768 18656 55820
rect 17776 55743 17828 55752
rect 17776 55709 17785 55743
rect 17785 55709 17819 55743
rect 17819 55709 17828 55743
rect 17776 55700 17828 55709
rect 18328 55743 18380 55752
rect 18328 55709 18337 55743
rect 18337 55709 18371 55743
rect 18371 55709 18380 55743
rect 18328 55700 18380 55709
rect 19524 55768 19576 55820
rect 20536 55768 20588 55820
rect 22100 55768 22152 55820
rect 24768 55768 24820 55820
rect 26976 55768 27028 55820
rect 30104 55811 30156 55820
rect 30104 55777 30113 55811
rect 30113 55777 30147 55811
rect 30147 55777 30156 55811
rect 30104 55768 30156 55777
rect 52920 55904 52972 55956
rect 55312 55904 55364 55956
rect 19708 55743 19760 55752
rect 19708 55709 19717 55743
rect 19717 55709 19751 55743
rect 19751 55709 19760 55743
rect 19708 55700 19760 55709
rect 22008 55700 22060 55752
rect 23848 55700 23900 55752
rect 19616 55675 19668 55684
rect 19616 55641 19625 55675
rect 19625 55641 19659 55675
rect 19659 55641 19668 55675
rect 19616 55632 19668 55641
rect 15936 55607 15988 55616
rect 15936 55573 15945 55607
rect 15945 55573 15979 55607
rect 15979 55573 15988 55607
rect 15936 55564 15988 55573
rect 16764 55564 16816 55616
rect 16948 55607 17000 55616
rect 16948 55573 16957 55607
rect 16957 55573 16991 55607
rect 16991 55573 17000 55607
rect 16948 55564 17000 55573
rect 17224 55564 17276 55616
rect 20628 55564 20680 55616
rect 22376 55607 22428 55616
rect 22376 55573 22385 55607
rect 22385 55573 22419 55607
rect 22419 55573 22428 55607
rect 22376 55564 22428 55573
rect 22744 55675 22796 55684
rect 22744 55641 22753 55675
rect 22753 55641 22787 55675
rect 22787 55641 22796 55675
rect 22744 55632 22796 55641
rect 26240 55743 26292 55752
rect 26240 55709 26249 55743
rect 26249 55709 26283 55743
rect 26283 55709 26292 55743
rect 26240 55700 26292 55709
rect 28080 55743 28132 55752
rect 28080 55709 28089 55743
rect 28089 55709 28123 55743
rect 28123 55709 28132 55743
rect 28080 55700 28132 55709
rect 43444 55743 43496 55752
rect 43444 55709 43453 55743
rect 43453 55709 43487 55743
rect 43487 55709 43496 55743
rect 43444 55700 43496 55709
rect 43904 55700 43956 55752
rect 44364 55743 44416 55752
rect 44364 55709 44373 55743
rect 44373 55709 44407 55743
rect 44407 55709 44416 55743
rect 44364 55700 44416 55709
rect 44916 55700 44968 55752
rect 45560 55743 45612 55752
rect 45560 55709 45569 55743
rect 45569 55709 45603 55743
rect 45603 55709 45612 55743
rect 45560 55700 45612 55709
rect 23020 55564 23072 55616
rect 23112 55564 23164 55616
rect 26424 55632 26476 55684
rect 27804 55632 27856 55684
rect 36176 55632 36228 55684
rect 38016 55675 38068 55684
rect 38016 55641 38025 55675
rect 38025 55641 38059 55675
rect 38059 55641 38068 55675
rect 38016 55632 38068 55641
rect 44732 55632 44784 55684
rect 51632 55811 51684 55820
rect 51632 55777 51641 55811
rect 51641 55777 51675 55811
rect 51675 55777 51684 55811
rect 51632 55768 51684 55777
rect 51356 55743 51408 55752
rect 51356 55709 51365 55743
rect 51365 55709 51399 55743
rect 51399 55709 51408 55743
rect 51356 55700 51408 55709
rect 24492 55607 24544 55616
rect 24492 55573 24501 55607
rect 24501 55573 24535 55607
rect 24535 55573 24544 55607
rect 24492 55564 24544 55573
rect 28448 55564 28500 55616
rect 29552 55564 29604 55616
rect 33416 55564 33468 55616
rect 35532 55564 35584 55616
rect 43260 55607 43312 55616
rect 43260 55573 43269 55607
rect 43269 55573 43303 55607
rect 43303 55573 43312 55607
rect 43260 55564 43312 55573
rect 44548 55607 44600 55616
rect 44548 55573 44557 55607
rect 44557 55573 44591 55607
rect 44591 55573 44600 55607
rect 44548 55564 44600 55573
rect 44640 55607 44692 55616
rect 44640 55573 44649 55607
rect 44649 55573 44683 55607
rect 44683 55573 44692 55607
rect 44640 55564 44692 55573
rect 49608 55564 49660 55616
rect 51540 55564 51592 55616
rect 52644 55564 52696 55616
rect 3010 55462 3062 55514
rect 3074 55462 3126 55514
rect 3138 55462 3190 55514
rect 3202 55462 3254 55514
rect 3266 55462 3318 55514
rect 33730 55462 33782 55514
rect 33794 55462 33846 55514
rect 33858 55462 33910 55514
rect 33922 55462 33974 55514
rect 33986 55462 34038 55514
rect 19708 55360 19760 55412
rect 19800 55360 19852 55412
rect 16856 55292 16908 55344
rect 16764 55224 16816 55276
rect 19616 55292 19668 55344
rect 16948 55199 17000 55208
rect 16948 55165 16957 55199
rect 16957 55165 16991 55199
rect 16991 55165 17000 55199
rect 16948 55156 17000 55165
rect 17500 55267 17552 55276
rect 17500 55233 17509 55267
rect 17509 55233 17543 55267
rect 17543 55233 17552 55267
rect 17500 55224 17552 55233
rect 22100 55360 22152 55412
rect 22468 55360 22520 55412
rect 20904 55292 20956 55344
rect 22008 55292 22060 55344
rect 23112 55292 23164 55344
rect 24492 55292 24544 55344
rect 22100 55224 22152 55276
rect 22284 55224 22336 55276
rect 22836 55224 22888 55276
rect 23020 55224 23072 55276
rect 17960 55156 18012 55208
rect 19892 55156 19944 55208
rect 21824 55199 21876 55208
rect 21824 55165 21833 55199
rect 21833 55165 21867 55199
rect 21867 55165 21876 55199
rect 21824 55156 21876 55165
rect 26332 55360 26384 55412
rect 27068 55360 27120 55412
rect 25044 55335 25096 55344
rect 25044 55301 25053 55335
rect 25053 55301 25087 55335
rect 25087 55301 25096 55335
rect 25044 55292 25096 55301
rect 26424 55292 26476 55344
rect 27804 55292 27856 55344
rect 24768 55199 24820 55208
rect 24768 55165 24777 55199
rect 24777 55165 24811 55199
rect 24811 55165 24820 55199
rect 24768 55156 24820 55165
rect 19984 55020 20036 55072
rect 23296 55020 23348 55072
rect 26516 55224 26568 55276
rect 28448 55335 28500 55344
rect 28448 55301 28457 55335
rect 28457 55301 28491 55335
rect 28491 55301 28500 55335
rect 28448 55292 28500 55301
rect 29552 55224 29604 55276
rect 32036 55360 32088 55412
rect 32404 55335 32456 55344
rect 32404 55301 32413 55335
rect 32413 55301 32447 55335
rect 32447 55301 32456 55335
rect 32404 55292 32456 55301
rect 33416 55292 33468 55344
rect 35900 55360 35952 55412
rect 37924 55360 37976 55412
rect 38476 55360 38528 55412
rect 35532 55292 35584 55344
rect 37280 55292 37332 55344
rect 40224 55360 40276 55412
rect 41604 55403 41656 55412
rect 41604 55369 41613 55403
rect 41613 55369 41647 55403
rect 41647 55369 41656 55403
rect 41604 55360 41656 55369
rect 43260 55335 43312 55344
rect 43260 55301 43269 55335
rect 43269 55301 43303 55335
rect 43303 55301 43312 55335
rect 43260 55292 43312 55301
rect 37924 55224 37976 55276
rect 34796 55156 34848 55208
rect 34244 55020 34296 55072
rect 38384 55156 38436 55208
rect 40132 55199 40184 55208
rect 40132 55165 40141 55199
rect 40141 55165 40175 55199
rect 40175 55165 40184 55199
rect 40132 55156 40184 55165
rect 42984 55199 43036 55208
rect 42984 55165 42993 55199
rect 42993 55165 43027 55199
rect 43027 55165 43036 55199
rect 42984 55156 43036 55165
rect 44272 55156 44324 55208
rect 44732 55403 44784 55412
rect 44732 55369 44741 55403
rect 44741 55369 44775 55403
rect 44775 55369 44784 55403
rect 44732 55360 44784 55369
rect 46756 55360 46808 55412
rect 48596 55292 48648 55344
rect 44548 55156 44600 55208
rect 45192 55156 45244 55208
rect 46756 55224 46808 55276
rect 48780 55292 48832 55344
rect 49608 55292 49660 55344
rect 51356 55360 51408 55412
rect 51080 55335 51132 55344
rect 51080 55301 51089 55335
rect 51089 55301 51123 55335
rect 51123 55301 51132 55335
rect 51080 55292 51132 55301
rect 51540 55292 51592 55344
rect 55220 55360 55272 55412
rect 52920 55292 52972 55344
rect 53472 55292 53524 55344
rect 46940 55156 46992 55208
rect 49792 55156 49844 55208
rect 51172 55156 51224 55208
rect 51724 55156 51776 55208
rect 39856 55088 39908 55140
rect 52552 55199 52604 55208
rect 52552 55165 52561 55199
rect 52561 55165 52595 55199
rect 52595 55165 52604 55199
rect 52552 55156 52604 55165
rect 38016 55020 38068 55072
rect 38660 55020 38712 55072
rect 2350 54918 2402 54970
rect 2414 54918 2466 54970
rect 2478 54918 2530 54970
rect 2542 54918 2594 54970
rect 2606 54918 2658 54970
rect 33070 54918 33122 54970
rect 33134 54918 33186 54970
rect 33198 54918 33250 54970
rect 33262 54918 33314 54970
rect 33326 54918 33378 54970
rect 20444 54816 20496 54868
rect 19340 54748 19392 54800
rect 22468 54723 22520 54732
rect 22468 54689 22477 54723
rect 22477 54689 22511 54723
rect 22511 54689 22520 54723
rect 22468 54680 22520 54689
rect 23296 54816 23348 54868
rect 30104 54816 30156 54868
rect 36268 54859 36320 54868
rect 36268 54825 36277 54859
rect 36277 54825 36311 54859
rect 36311 54825 36320 54859
rect 36268 54816 36320 54825
rect 39856 54816 39908 54868
rect 26240 54791 26292 54800
rect 26240 54757 26249 54791
rect 26249 54757 26283 54791
rect 26283 54757 26292 54791
rect 26240 54748 26292 54757
rect 27896 54723 27948 54732
rect 27896 54689 27905 54723
rect 27905 54689 27939 54723
rect 27939 54689 27948 54723
rect 27896 54680 27948 54689
rect 37740 54723 37792 54732
rect 37740 54689 37749 54723
rect 37749 54689 37783 54723
rect 37783 54689 37792 54723
rect 37740 54680 37792 54689
rect 38016 54723 38068 54732
rect 38016 54689 38025 54723
rect 38025 54689 38059 54723
rect 38059 54689 38068 54723
rect 38016 54680 38068 54689
rect 43904 54816 43956 54868
rect 53012 54816 53064 54868
rect 42984 54680 43036 54732
rect 46756 54723 46808 54732
rect 46756 54689 46765 54723
rect 46765 54689 46799 54723
rect 46799 54689 46808 54723
rect 46756 54680 46808 54689
rect 51356 54723 51408 54732
rect 51356 54689 51365 54723
rect 51365 54689 51399 54723
rect 51399 54689 51408 54723
rect 51356 54680 51408 54689
rect 52000 54680 52052 54732
rect 52644 54680 52696 54732
rect 23848 54612 23900 54664
rect 29552 54612 29604 54664
rect 44272 54612 44324 54664
rect 44824 54612 44876 54664
rect 45192 54612 45244 54664
rect 22008 54544 22060 54596
rect 15936 54476 15988 54528
rect 27804 54476 27856 54528
rect 36176 54544 36228 54596
rect 37280 54544 37332 54596
rect 41972 54587 42024 54596
rect 41972 54553 41981 54587
rect 41981 54553 42015 54587
rect 42015 54553 42024 54587
rect 41972 54544 42024 54553
rect 53472 54612 53524 54664
rect 58256 54612 58308 54664
rect 3010 54374 3062 54426
rect 3074 54374 3126 54426
rect 3138 54374 3190 54426
rect 3202 54374 3254 54426
rect 3266 54374 3318 54426
rect 33730 54374 33782 54426
rect 33794 54374 33846 54426
rect 33858 54374 33910 54426
rect 33922 54374 33974 54426
rect 33986 54374 34038 54426
rect 19616 54272 19668 54324
rect 21088 54204 21140 54256
rect 22008 54204 22060 54256
rect 46756 54272 46808 54324
rect 44640 54204 44692 54256
rect 44824 54204 44876 54256
rect 20812 54068 20864 54120
rect 22468 54068 22520 54120
rect 45836 54111 45888 54120
rect 45836 54077 45845 54111
rect 45845 54077 45879 54111
rect 45879 54077 45888 54111
rect 45836 54068 45888 54077
rect 16212 53932 16264 53984
rect 2350 53830 2402 53882
rect 2414 53830 2466 53882
rect 2478 53830 2530 53882
rect 2542 53830 2594 53882
rect 2606 53830 2658 53882
rect 33070 53830 33122 53882
rect 33134 53830 33186 53882
rect 33198 53830 33250 53882
rect 33262 53830 33314 53882
rect 33326 53830 33378 53882
rect 17776 53728 17828 53780
rect 26516 53771 26568 53780
rect 26516 53737 26525 53771
rect 26525 53737 26559 53771
rect 26559 53737 26568 53771
rect 26516 53728 26568 53737
rect 22468 53635 22520 53644
rect 22468 53601 22477 53635
rect 22477 53601 22511 53635
rect 22511 53601 22520 53635
rect 22468 53592 22520 53601
rect 21088 53524 21140 53576
rect 27804 53567 27856 53576
rect 27804 53533 27813 53567
rect 27813 53533 27847 53567
rect 27847 53533 27856 53567
rect 27804 53524 27856 53533
rect 22560 53456 22612 53508
rect 3010 53286 3062 53338
rect 3074 53286 3126 53338
rect 3138 53286 3190 53338
rect 3202 53286 3254 53338
rect 3266 53286 3318 53338
rect 33730 53286 33782 53338
rect 33794 53286 33846 53338
rect 33858 53286 33910 53338
rect 33922 53286 33974 53338
rect 33986 53286 34038 53338
rect 19432 53184 19484 53236
rect 21088 53116 21140 53168
rect 22468 53048 22520 53100
rect 20628 52980 20680 53032
rect 2350 52742 2402 52794
rect 2414 52742 2466 52794
rect 2478 52742 2530 52794
rect 2542 52742 2594 52794
rect 2606 52742 2658 52794
rect 33070 52742 33122 52794
rect 33134 52742 33186 52794
rect 33198 52742 33250 52794
rect 33262 52742 33314 52794
rect 33326 52742 33378 52794
rect 3010 52198 3062 52250
rect 3074 52198 3126 52250
rect 3138 52198 3190 52250
rect 3202 52198 3254 52250
rect 3266 52198 3318 52250
rect 33730 52198 33782 52250
rect 33794 52198 33846 52250
rect 33858 52198 33910 52250
rect 33922 52198 33974 52250
rect 33986 52198 34038 52250
rect 2350 51654 2402 51706
rect 2414 51654 2466 51706
rect 2478 51654 2530 51706
rect 2542 51654 2594 51706
rect 2606 51654 2658 51706
rect 33070 51654 33122 51706
rect 33134 51654 33186 51706
rect 33198 51654 33250 51706
rect 33262 51654 33314 51706
rect 33326 51654 33378 51706
rect 3010 51110 3062 51162
rect 3074 51110 3126 51162
rect 3138 51110 3190 51162
rect 3202 51110 3254 51162
rect 3266 51110 3318 51162
rect 33730 51110 33782 51162
rect 33794 51110 33846 51162
rect 33858 51110 33910 51162
rect 33922 51110 33974 51162
rect 33986 51110 34038 51162
rect 2350 50566 2402 50618
rect 2414 50566 2466 50618
rect 2478 50566 2530 50618
rect 2542 50566 2594 50618
rect 2606 50566 2658 50618
rect 33070 50566 33122 50618
rect 33134 50566 33186 50618
rect 33198 50566 33250 50618
rect 33262 50566 33314 50618
rect 33326 50566 33378 50618
rect 3010 50022 3062 50074
rect 3074 50022 3126 50074
rect 3138 50022 3190 50074
rect 3202 50022 3254 50074
rect 3266 50022 3318 50074
rect 33730 50022 33782 50074
rect 33794 50022 33846 50074
rect 33858 50022 33910 50074
rect 33922 50022 33974 50074
rect 33986 50022 34038 50074
rect 2350 49478 2402 49530
rect 2414 49478 2466 49530
rect 2478 49478 2530 49530
rect 2542 49478 2594 49530
rect 2606 49478 2658 49530
rect 33070 49478 33122 49530
rect 33134 49478 33186 49530
rect 33198 49478 33250 49530
rect 33262 49478 33314 49530
rect 33326 49478 33378 49530
rect 3010 48934 3062 48986
rect 3074 48934 3126 48986
rect 3138 48934 3190 48986
rect 3202 48934 3254 48986
rect 3266 48934 3318 48986
rect 33730 48934 33782 48986
rect 33794 48934 33846 48986
rect 33858 48934 33910 48986
rect 33922 48934 33974 48986
rect 33986 48934 34038 48986
rect 2350 48390 2402 48442
rect 2414 48390 2466 48442
rect 2478 48390 2530 48442
rect 2542 48390 2594 48442
rect 2606 48390 2658 48442
rect 33070 48390 33122 48442
rect 33134 48390 33186 48442
rect 33198 48390 33250 48442
rect 33262 48390 33314 48442
rect 33326 48390 33378 48442
rect 3010 47846 3062 47898
rect 3074 47846 3126 47898
rect 3138 47846 3190 47898
rect 3202 47846 3254 47898
rect 3266 47846 3318 47898
rect 33730 47846 33782 47898
rect 33794 47846 33846 47898
rect 33858 47846 33910 47898
rect 33922 47846 33974 47898
rect 33986 47846 34038 47898
rect 2350 47302 2402 47354
rect 2414 47302 2466 47354
rect 2478 47302 2530 47354
rect 2542 47302 2594 47354
rect 2606 47302 2658 47354
rect 33070 47302 33122 47354
rect 33134 47302 33186 47354
rect 33198 47302 33250 47354
rect 33262 47302 33314 47354
rect 33326 47302 33378 47354
rect 3010 46758 3062 46810
rect 3074 46758 3126 46810
rect 3138 46758 3190 46810
rect 3202 46758 3254 46810
rect 3266 46758 3318 46810
rect 33730 46758 33782 46810
rect 33794 46758 33846 46810
rect 33858 46758 33910 46810
rect 33922 46758 33974 46810
rect 33986 46758 34038 46810
rect 2350 46214 2402 46266
rect 2414 46214 2466 46266
rect 2478 46214 2530 46266
rect 2542 46214 2594 46266
rect 2606 46214 2658 46266
rect 33070 46214 33122 46266
rect 33134 46214 33186 46266
rect 33198 46214 33250 46266
rect 33262 46214 33314 46266
rect 33326 46214 33378 46266
rect 3010 45670 3062 45722
rect 3074 45670 3126 45722
rect 3138 45670 3190 45722
rect 3202 45670 3254 45722
rect 3266 45670 3318 45722
rect 33730 45670 33782 45722
rect 33794 45670 33846 45722
rect 33858 45670 33910 45722
rect 33922 45670 33974 45722
rect 33986 45670 34038 45722
rect 2350 45126 2402 45178
rect 2414 45126 2466 45178
rect 2478 45126 2530 45178
rect 2542 45126 2594 45178
rect 2606 45126 2658 45178
rect 33070 45126 33122 45178
rect 33134 45126 33186 45178
rect 33198 45126 33250 45178
rect 33262 45126 33314 45178
rect 33326 45126 33378 45178
rect 58256 44931 58308 44940
rect 58256 44897 58265 44931
rect 58265 44897 58299 44931
rect 58299 44897 58308 44931
rect 58256 44888 58308 44897
rect 58532 44863 58584 44872
rect 58532 44829 58541 44863
rect 58541 44829 58575 44863
rect 58575 44829 58584 44863
rect 58532 44820 58584 44829
rect 3010 44582 3062 44634
rect 3074 44582 3126 44634
rect 3138 44582 3190 44634
rect 3202 44582 3254 44634
rect 3266 44582 3318 44634
rect 33730 44582 33782 44634
rect 33794 44582 33846 44634
rect 33858 44582 33910 44634
rect 33922 44582 33974 44634
rect 33986 44582 34038 44634
rect 2350 44038 2402 44090
rect 2414 44038 2466 44090
rect 2478 44038 2530 44090
rect 2542 44038 2594 44090
rect 2606 44038 2658 44090
rect 33070 44038 33122 44090
rect 33134 44038 33186 44090
rect 33198 44038 33250 44090
rect 33262 44038 33314 44090
rect 33326 44038 33378 44090
rect 3010 43494 3062 43546
rect 3074 43494 3126 43546
rect 3138 43494 3190 43546
rect 3202 43494 3254 43546
rect 3266 43494 3318 43546
rect 33730 43494 33782 43546
rect 33794 43494 33846 43546
rect 33858 43494 33910 43546
rect 33922 43494 33974 43546
rect 33986 43494 34038 43546
rect 2350 42950 2402 43002
rect 2414 42950 2466 43002
rect 2478 42950 2530 43002
rect 2542 42950 2594 43002
rect 2606 42950 2658 43002
rect 33070 42950 33122 43002
rect 33134 42950 33186 43002
rect 33198 42950 33250 43002
rect 33262 42950 33314 43002
rect 33326 42950 33378 43002
rect 3010 42406 3062 42458
rect 3074 42406 3126 42458
rect 3138 42406 3190 42458
rect 3202 42406 3254 42458
rect 3266 42406 3318 42458
rect 33730 42406 33782 42458
rect 33794 42406 33846 42458
rect 33858 42406 33910 42458
rect 33922 42406 33974 42458
rect 33986 42406 34038 42458
rect 2350 41862 2402 41914
rect 2414 41862 2466 41914
rect 2478 41862 2530 41914
rect 2542 41862 2594 41914
rect 2606 41862 2658 41914
rect 33070 41862 33122 41914
rect 33134 41862 33186 41914
rect 33198 41862 33250 41914
rect 33262 41862 33314 41914
rect 33326 41862 33378 41914
rect 3010 41318 3062 41370
rect 3074 41318 3126 41370
rect 3138 41318 3190 41370
rect 3202 41318 3254 41370
rect 3266 41318 3318 41370
rect 33730 41318 33782 41370
rect 33794 41318 33846 41370
rect 33858 41318 33910 41370
rect 33922 41318 33974 41370
rect 33986 41318 34038 41370
rect 2350 40774 2402 40826
rect 2414 40774 2466 40826
rect 2478 40774 2530 40826
rect 2542 40774 2594 40826
rect 2606 40774 2658 40826
rect 33070 40774 33122 40826
rect 33134 40774 33186 40826
rect 33198 40774 33250 40826
rect 33262 40774 33314 40826
rect 33326 40774 33378 40826
rect 3010 40230 3062 40282
rect 3074 40230 3126 40282
rect 3138 40230 3190 40282
rect 3202 40230 3254 40282
rect 3266 40230 3318 40282
rect 33730 40230 33782 40282
rect 33794 40230 33846 40282
rect 33858 40230 33910 40282
rect 33922 40230 33974 40282
rect 33986 40230 34038 40282
rect 2350 39686 2402 39738
rect 2414 39686 2466 39738
rect 2478 39686 2530 39738
rect 2542 39686 2594 39738
rect 2606 39686 2658 39738
rect 33070 39686 33122 39738
rect 33134 39686 33186 39738
rect 33198 39686 33250 39738
rect 33262 39686 33314 39738
rect 33326 39686 33378 39738
rect 3010 39142 3062 39194
rect 3074 39142 3126 39194
rect 3138 39142 3190 39194
rect 3202 39142 3254 39194
rect 3266 39142 3318 39194
rect 33730 39142 33782 39194
rect 33794 39142 33846 39194
rect 33858 39142 33910 39194
rect 33922 39142 33974 39194
rect 33986 39142 34038 39194
rect 2350 38598 2402 38650
rect 2414 38598 2466 38650
rect 2478 38598 2530 38650
rect 2542 38598 2594 38650
rect 2606 38598 2658 38650
rect 33070 38598 33122 38650
rect 33134 38598 33186 38650
rect 33198 38598 33250 38650
rect 33262 38598 33314 38650
rect 33326 38598 33378 38650
rect 3010 38054 3062 38106
rect 3074 38054 3126 38106
rect 3138 38054 3190 38106
rect 3202 38054 3254 38106
rect 3266 38054 3318 38106
rect 33730 38054 33782 38106
rect 33794 38054 33846 38106
rect 33858 38054 33910 38106
rect 33922 38054 33974 38106
rect 33986 38054 34038 38106
rect 2350 37510 2402 37562
rect 2414 37510 2466 37562
rect 2478 37510 2530 37562
rect 2542 37510 2594 37562
rect 2606 37510 2658 37562
rect 33070 37510 33122 37562
rect 33134 37510 33186 37562
rect 33198 37510 33250 37562
rect 33262 37510 33314 37562
rect 33326 37510 33378 37562
rect 3010 36966 3062 37018
rect 3074 36966 3126 37018
rect 3138 36966 3190 37018
rect 3202 36966 3254 37018
rect 3266 36966 3318 37018
rect 33730 36966 33782 37018
rect 33794 36966 33846 37018
rect 33858 36966 33910 37018
rect 33922 36966 33974 37018
rect 33986 36966 34038 37018
rect 2350 36422 2402 36474
rect 2414 36422 2466 36474
rect 2478 36422 2530 36474
rect 2542 36422 2594 36474
rect 2606 36422 2658 36474
rect 33070 36422 33122 36474
rect 33134 36422 33186 36474
rect 33198 36422 33250 36474
rect 33262 36422 33314 36474
rect 33326 36422 33378 36474
rect 3010 35878 3062 35930
rect 3074 35878 3126 35930
rect 3138 35878 3190 35930
rect 3202 35878 3254 35930
rect 3266 35878 3318 35930
rect 33730 35878 33782 35930
rect 33794 35878 33846 35930
rect 33858 35878 33910 35930
rect 33922 35878 33974 35930
rect 33986 35878 34038 35930
rect 2350 35334 2402 35386
rect 2414 35334 2466 35386
rect 2478 35334 2530 35386
rect 2542 35334 2594 35386
rect 2606 35334 2658 35386
rect 33070 35334 33122 35386
rect 33134 35334 33186 35386
rect 33198 35334 33250 35386
rect 33262 35334 33314 35386
rect 33326 35334 33378 35386
rect 3010 34790 3062 34842
rect 3074 34790 3126 34842
rect 3138 34790 3190 34842
rect 3202 34790 3254 34842
rect 3266 34790 3318 34842
rect 33730 34790 33782 34842
rect 33794 34790 33846 34842
rect 33858 34790 33910 34842
rect 33922 34790 33974 34842
rect 33986 34790 34038 34842
rect 2350 34246 2402 34298
rect 2414 34246 2466 34298
rect 2478 34246 2530 34298
rect 2542 34246 2594 34298
rect 2606 34246 2658 34298
rect 33070 34246 33122 34298
rect 33134 34246 33186 34298
rect 33198 34246 33250 34298
rect 33262 34246 33314 34298
rect 33326 34246 33378 34298
rect 3010 33702 3062 33754
rect 3074 33702 3126 33754
rect 3138 33702 3190 33754
rect 3202 33702 3254 33754
rect 3266 33702 3318 33754
rect 33730 33702 33782 33754
rect 33794 33702 33846 33754
rect 33858 33702 33910 33754
rect 33922 33702 33974 33754
rect 33986 33702 34038 33754
rect 2350 33158 2402 33210
rect 2414 33158 2466 33210
rect 2478 33158 2530 33210
rect 2542 33158 2594 33210
rect 2606 33158 2658 33210
rect 33070 33158 33122 33210
rect 33134 33158 33186 33210
rect 33198 33158 33250 33210
rect 33262 33158 33314 33210
rect 33326 33158 33378 33210
rect 3010 32614 3062 32666
rect 3074 32614 3126 32666
rect 3138 32614 3190 32666
rect 3202 32614 3254 32666
rect 3266 32614 3318 32666
rect 33730 32614 33782 32666
rect 33794 32614 33846 32666
rect 33858 32614 33910 32666
rect 33922 32614 33974 32666
rect 33986 32614 34038 32666
rect 2350 32070 2402 32122
rect 2414 32070 2466 32122
rect 2478 32070 2530 32122
rect 2542 32070 2594 32122
rect 2606 32070 2658 32122
rect 33070 32070 33122 32122
rect 33134 32070 33186 32122
rect 33198 32070 33250 32122
rect 33262 32070 33314 32122
rect 33326 32070 33378 32122
rect 3010 31526 3062 31578
rect 3074 31526 3126 31578
rect 3138 31526 3190 31578
rect 3202 31526 3254 31578
rect 3266 31526 3318 31578
rect 33730 31526 33782 31578
rect 33794 31526 33846 31578
rect 33858 31526 33910 31578
rect 33922 31526 33974 31578
rect 33986 31526 34038 31578
rect 2350 30982 2402 31034
rect 2414 30982 2466 31034
rect 2478 30982 2530 31034
rect 2542 30982 2594 31034
rect 2606 30982 2658 31034
rect 33070 30982 33122 31034
rect 33134 30982 33186 31034
rect 33198 30982 33250 31034
rect 33262 30982 33314 31034
rect 33326 30982 33378 31034
rect 3010 30438 3062 30490
rect 3074 30438 3126 30490
rect 3138 30438 3190 30490
rect 3202 30438 3254 30490
rect 3266 30438 3318 30490
rect 33730 30438 33782 30490
rect 33794 30438 33846 30490
rect 33858 30438 33910 30490
rect 33922 30438 33974 30490
rect 33986 30438 34038 30490
rect 2350 29894 2402 29946
rect 2414 29894 2466 29946
rect 2478 29894 2530 29946
rect 2542 29894 2594 29946
rect 2606 29894 2658 29946
rect 33070 29894 33122 29946
rect 33134 29894 33186 29946
rect 33198 29894 33250 29946
rect 33262 29894 33314 29946
rect 33326 29894 33378 29946
rect 3010 29350 3062 29402
rect 3074 29350 3126 29402
rect 3138 29350 3190 29402
rect 3202 29350 3254 29402
rect 3266 29350 3318 29402
rect 33730 29350 33782 29402
rect 33794 29350 33846 29402
rect 33858 29350 33910 29402
rect 33922 29350 33974 29402
rect 33986 29350 34038 29402
rect 2350 28806 2402 28858
rect 2414 28806 2466 28858
rect 2478 28806 2530 28858
rect 2542 28806 2594 28858
rect 2606 28806 2658 28858
rect 33070 28806 33122 28858
rect 33134 28806 33186 28858
rect 33198 28806 33250 28858
rect 33262 28806 33314 28858
rect 33326 28806 33378 28858
rect 3010 28262 3062 28314
rect 3074 28262 3126 28314
rect 3138 28262 3190 28314
rect 3202 28262 3254 28314
rect 3266 28262 3318 28314
rect 33730 28262 33782 28314
rect 33794 28262 33846 28314
rect 33858 28262 33910 28314
rect 33922 28262 33974 28314
rect 33986 28262 34038 28314
rect 2350 27718 2402 27770
rect 2414 27718 2466 27770
rect 2478 27718 2530 27770
rect 2542 27718 2594 27770
rect 2606 27718 2658 27770
rect 33070 27718 33122 27770
rect 33134 27718 33186 27770
rect 33198 27718 33250 27770
rect 33262 27718 33314 27770
rect 33326 27718 33378 27770
rect 3010 27174 3062 27226
rect 3074 27174 3126 27226
rect 3138 27174 3190 27226
rect 3202 27174 3254 27226
rect 3266 27174 3318 27226
rect 33730 27174 33782 27226
rect 33794 27174 33846 27226
rect 33858 27174 33910 27226
rect 33922 27174 33974 27226
rect 33986 27174 34038 27226
rect 2350 26630 2402 26682
rect 2414 26630 2466 26682
rect 2478 26630 2530 26682
rect 2542 26630 2594 26682
rect 2606 26630 2658 26682
rect 33070 26630 33122 26682
rect 33134 26630 33186 26682
rect 33198 26630 33250 26682
rect 33262 26630 33314 26682
rect 33326 26630 33378 26682
rect 3010 26086 3062 26138
rect 3074 26086 3126 26138
rect 3138 26086 3190 26138
rect 3202 26086 3254 26138
rect 3266 26086 3318 26138
rect 33730 26086 33782 26138
rect 33794 26086 33846 26138
rect 33858 26086 33910 26138
rect 33922 26086 33974 26138
rect 33986 26086 34038 26138
rect 2350 25542 2402 25594
rect 2414 25542 2466 25594
rect 2478 25542 2530 25594
rect 2542 25542 2594 25594
rect 2606 25542 2658 25594
rect 33070 25542 33122 25594
rect 33134 25542 33186 25594
rect 33198 25542 33250 25594
rect 33262 25542 33314 25594
rect 33326 25542 33378 25594
rect 3010 24998 3062 25050
rect 3074 24998 3126 25050
rect 3138 24998 3190 25050
rect 3202 24998 3254 25050
rect 3266 24998 3318 25050
rect 33730 24998 33782 25050
rect 33794 24998 33846 25050
rect 33858 24998 33910 25050
rect 33922 24998 33974 25050
rect 33986 24998 34038 25050
rect 2350 24454 2402 24506
rect 2414 24454 2466 24506
rect 2478 24454 2530 24506
rect 2542 24454 2594 24506
rect 2606 24454 2658 24506
rect 33070 24454 33122 24506
rect 33134 24454 33186 24506
rect 33198 24454 33250 24506
rect 33262 24454 33314 24506
rect 33326 24454 33378 24506
rect 3010 23910 3062 23962
rect 3074 23910 3126 23962
rect 3138 23910 3190 23962
rect 3202 23910 3254 23962
rect 3266 23910 3318 23962
rect 33730 23910 33782 23962
rect 33794 23910 33846 23962
rect 33858 23910 33910 23962
rect 33922 23910 33974 23962
rect 33986 23910 34038 23962
rect 2350 23366 2402 23418
rect 2414 23366 2466 23418
rect 2478 23366 2530 23418
rect 2542 23366 2594 23418
rect 2606 23366 2658 23418
rect 33070 23366 33122 23418
rect 33134 23366 33186 23418
rect 33198 23366 33250 23418
rect 33262 23366 33314 23418
rect 33326 23366 33378 23418
rect 3010 22822 3062 22874
rect 3074 22822 3126 22874
rect 3138 22822 3190 22874
rect 3202 22822 3254 22874
rect 3266 22822 3318 22874
rect 33730 22822 33782 22874
rect 33794 22822 33846 22874
rect 33858 22822 33910 22874
rect 33922 22822 33974 22874
rect 33986 22822 34038 22874
rect 2350 22278 2402 22330
rect 2414 22278 2466 22330
rect 2478 22278 2530 22330
rect 2542 22278 2594 22330
rect 2606 22278 2658 22330
rect 33070 22278 33122 22330
rect 33134 22278 33186 22330
rect 33198 22278 33250 22330
rect 33262 22278 33314 22330
rect 33326 22278 33378 22330
rect 3010 21734 3062 21786
rect 3074 21734 3126 21786
rect 3138 21734 3190 21786
rect 3202 21734 3254 21786
rect 3266 21734 3318 21786
rect 33730 21734 33782 21786
rect 33794 21734 33846 21786
rect 33858 21734 33910 21786
rect 33922 21734 33974 21786
rect 33986 21734 34038 21786
rect 2350 21190 2402 21242
rect 2414 21190 2466 21242
rect 2478 21190 2530 21242
rect 2542 21190 2594 21242
rect 2606 21190 2658 21242
rect 33070 21190 33122 21242
rect 33134 21190 33186 21242
rect 33198 21190 33250 21242
rect 33262 21190 33314 21242
rect 33326 21190 33378 21242
rect 3010 20646 3062 20698
rect 3074 20646 3126 20698
rect 3138 20646 3190 20698
rect 3202 20646 3254 20698
rect 3266 20646 3318 20698
rect 33730 20646 33782 20698
rect 33794 20646 33846 20698
rect 33858 20646 33910 20698
rect 33922 20646 33974 20698
rect 33986 20646 34038 20698
rect 2350 20102 2402 20154
rect 2414 20102 2466 20154
rect 2478 20102 2530 20154
rect 2542 20102 2594 20154
rect 2606 20102 2658 20154
rect 33070 20102 33122 20154
rect 33134 20102 33186 20154
rect 33198 20102 33250 20154
rect 33262 20102 33314 20154
rect 33326 20102 33378 20154
rect 3010 19558 3062 19610
rect 3074 19558 3126 19610
rect 3138 19558 3190 19610
rect 3202 19558 3254 19610
rect 3266 19558 3318 19610
rect 33730 19558 33782 19610
rect 33794 19558 33846 19610
rect 33858 19558 33910 19610
rect 33922 19558 33974 19610
rect 33986 19558 34038 19610
rect 2350 19014 2402 19066
rect 2414 19014 2466 19066
rect 2478 19014 2530 19066
rect 2542 19014 2594 19066
rect 2606 19014 2658 19066
rect 33070 19014 33122 19066
rect 33134 19014 33186 19066
rect 33198 19014 33250 19066
rect 33262 19014 33314 19066
rect 33326 19014 33378 19066
rect 3010 18470 3062 18522
rect 3074 18470 3126 18522
rect 3138 18470 3190 18522
rect 3202 18470 3254 18522
rect 3266 18470 3318 18522
rect 33730 18470 33782 18522
rect 33794 18470 33846 18522
rect 33858 18470 33910 18522
rect 33922 18470 33974 18522
rect 33986 18470 34038 18522
rect 2350 17926 2402 17978
rect 2414 17926 2466 17978
rect 2478 17926 2530 17978
rect 2542 17926 2594 17978
rect 2606 17926 2658 17978
rect 33070 17926 33122 17978
rect 33134 17926 33186 17978
rect 33198 17926 33250 17978
rect 33262 17926 33314 17978
rect 33326 17926 33378 17978
rect 3010 17382 3062 17434
rect 3074 17382 3126 17434
rect 3138 17382 3190 17434
rect 3202 17382 3254 17434
rect 3266 17382 3318 17434
rect 33730 17382 33782 17434
rect 33794 17382 33846 17434
rect 33858 17382 33910 17434
rect 33922 17382 33974 17434
rect 33986 17382 34038 17434
rect 2350 16838 2402 16890
rect 2414 16838 2466 16890
rect 2478 16838 2530 16890
rect 2542 16838 2594 16890
rect 2606 16838 2658 16890
rect 33070 16838 33122 16890
rect 33134 16838 33186 16890
rect 33198 16838 33250 16890
rect 33262 16838 33314 16890
rect 33326 16838 33378 16890
rect 3010 16294 3062 16346
rect 3074 16294 3126 16346
rect 3138 16294 3190 16346
rect 3202 16294 3254 16346
rect 3266 16294 3318 16346
rect 33730 16294 33782 16346
rect 33794 16294 33846 16346
rect 33858 16294 33910 16346
rect 33922 16294 33974 16346
rect 33986 16294 34038 16346
rect 2350 15750 2402 15802
rect 2414 15750 2466 15802
rect 2478 15750 2530 15802
rect 2542 15750 2594 15802
rect 2606 15750 2658 15802
rect 33070 15750 33122 15802
rect 33134 15750 33186 15802
rect 33198 15750 33250 15802
rect 33262 15750 33314 15802
rect 33326 15750 33378 15802
rect 3010 15206 3062 15258
rect 3074 15206 3126 15258
rect 3138 15206 3190 15258
rect 3202 15206 3254 15258
rect 3266 15206 3318 15258
rect 33730 15206 33782 15258
rect 33794 15206 33846 15258
rect 33858 15206 33910 15258
rect 33922 15206 33974 15258
rect 33986 15206 34038 15258
rect 38016 15104 38068 15156
rect 56508 15104 56560 15156
rect 2350 14662 2402 14714
rect 2414 14662 2466 14714
rect 2478 14662 2530 14714
rect 2542 14662 2594 14714
rect 2606 14662 2658 14714
rect 33070 14662 33122 14714
rect 33134 14662 33186 14714
rect 33198 14662 33250 14714
rect 33262 14662 33314 14714
rect 33326 14662 33378 14714
rect 3010 14118 3062 14170
rect 3074 14118 3126 14170
rect 3138 14118 3190 14170
rect 3202 14118 3254 14170
rect 3266 14118 3318 14170
rect 33730 14118 33782 14170
rect 33794 14118 33846 14170
rect 33858 14118 33910 14170
rect 33922 14118 33974 14170
rect 33986 14118 34038 14170
rect 2350 13574 2402 13626
rect 2414 13574 2466 13626
rect 2478 13574 2530 13626
rect 2542 13574 2594 13626
rect 2606 13574 2658 13626
rect 33070 13574 33122 13626
rect 33134 13574 33186 13626
rect 33198 13574 33250 13626
rect 33262 13574 33314 13626
rect 33326 13574 33378 13626
rect 3010 13030 3062 13082
rect 3074 13030 3126 13082
rect 3138 13030 3190 13082
rect 3202 13030 3254 13082
rect 3266 13030 3318 13082
rect 33730 13030 33782 13082
rect 33794 13030 33846 13082
rect 33858 13030 33910 13082
rect 33922 13030 33974 13082
rect 33986 13030 34038 13082
rect 2350 12486 2402 12538
rect 2414 12486 2466 12538
rect 2478 12486 2530 12538
rect 2542 12486 2594 12538
rect 2606 12486 2658 12538
rect 33070 12486 33122 12538
rect 33134 12486 33186 12538
rect 33198 12486 33250 12538
rect 33262 12486 33314 12538
rect 33326 12486 33378 12538
rect 3010 11942 3062 11994
rect 3074 11942 3126 11994
rect 3138 11942 3190 11994
rect 3202 11942 3254 11994
rect 3266 11942 3318 11994
rect 33730 11942 33782 11994
rect 33794 11942 33846 11994
rect 33858 11942 33910 11994
rect 33922 11942 33974 11994
rect 33986 11942 34038 11994
rect 2350 11398 2402 11450
rect 2414 11398 2466 11450
rect 2478 11398 2530 11450
rect 2542 11398 2594 11450
rect 2606 11398 2658 11450
rect 33070 11398 33122 11450
rect 33134 11398 33186 11450
rect 33198 11398 33250 11450
rect 33262 11398 33314 11450
rect 33326 11398 33378 11450
rect 3010 10854 3062 10906
rect 3074 10854 3126 10906
rect 3138 10854 3190 10906
rect 3202 10854 3254 10906
rect 3266 10854 3318 10906
rect 33730 10854 33782 10906
rect 33794 10854 33846 10906
rect 33858 10854 33910 10906
rect 33922 10854 33974 10906
rect 33986 10854 34038 10906
rect 2350 10310 2402 10362
rect 2414 10310 2466 10362
rect 2478 10310 2530 10362
rect 2542 10310 2594 10362
rect 2606 10310 2658 10362
rect 33070 10310 33122 10362
rect 33134 10310 33186 10362
rect 33198 10310 33250 10362
rect 33262 10310 33314 10362
rect 33326 10310 33378 10362
rect 3010 9766 3062 9818
rect 3074 9766 3126 9818
rect 3138 9766 3190 9818
rect 3202 9766 3254 9818
rect 3266 9766 3318 9818
rect 33730 9766 33782 9818
rect 33794 9766 33846 9818
rect 33858 9766 33910 9818
rect 33922 9766 33974 9818
rect 33986 9766 34038 9818
rect 2350 9222 2402 9274
rect 2414 9222 2466 9274
rect 2478 9222 2530 9274
rect 2542 9222 2594 9274
rect 2606 9222 2658 9274
rect 33070 9222 33122 9274
rect 33134 9222 33186 9274
rect 33198 9222 33250 9274
rect 33262 9222 33314 9274
rect 33326 9222 33378 9274
rect 3010 8678 3062 8730
rect 3074 8678 3126 8730
rect 3138 8678 3190 8730
rect 3202 8678 3254 8730
rect 3266 8678 3318 8730
rect 33730 8678 33782 8730
rect 33794 8678 33846 8730
rect 33858 8678 33910 8730
rect 33922 8678 33974 8730
rect 33986 8678 34038 8730
rect 2350 8134 2402 8186
rect 2414 8134 2466 8186
rect 2478 8134 2530 8186
rect 2542 8134 2594 8186
rect 2606 8134 2658 8186
rect 33070 8134 33122 8186
rect 33134 8134 33186 8186
rect 33198 8134 33250 8186
rect 33262 8134 33314 8186
rect 33326 8134 33378 8186
rect 3010 7590 3062 7642
rect 3074 7590 3126 7642
rect 3138 7590 3190 7642
rect 3202 7590 3254 7642
rect 3266 7590 3318 7642
rect 33730 7590 33782 7642
rect 33794 7590 33846 7642
rect 33858 7590 33910 7642
rect 33922 7590 33974 7642
rect 33986 7590 34038 7642
rect 2350 7046 2402 7098
rect 2414 7046 2466 7098
rect 2478 7046 2530 7098
rect 2542 7046 2594 7098
rect 2606 7046 2658 7098
rect 33070 7046 33122 7098
rect 33134 7046 33186 7098
rect 33198 7046 33250 7098
rect 33262 7046 33314 7098
rect 33326 7046 33378 7098
rect 3010 6502 3062 6554
rect 3074 6502 3126 6554
rect 3138 6502 3190 6554
rect 3202 6502 3254 6554
rect 3266 6502 3318 6554
rect 33730 6502 33782 6554
rect 33794 6502 33846 6554
rect 33858 6502 33910 6554
rect 33922 6502 33974 6554
rect 33986 6502 34038 6554
rect 2350 5958 2402 6010
rect 2414 5958 2466 6010
rect 2478 5958 2530 6010
rect 2542 5958 2594 6010
rect 2606 5958 2658 6010
rect 33070 5958 33122 6010
rect 33134 5958 33186 6010
rect 33198 5958 33250 6010
rect 33262 5958 33314 6010
rect 33326 5958 33378 6010
rect 3010 5414 3062 5466
rect 3074 5414 3126 5466
rect 3138 5414 3190 5466
rect 3202 5414 3254 5466
rect 3266 5414 3318 5466
rect 33730 5414 33782 5466
rect 33794 5414 33846 5466
rect 33858 5414 33910 5466
rect 33922 5414 33974 5466
rect 33986 5414 34038 5466
rect 2350 4870 2402 4922
rect 2414 4870 2466 4922
rect 2478 4870 2530 4922
rect 2542 4870 2594 4922
rect 2606 4870 2658 4922
rect 33070 4870 33122 4922
rect 33134 4870 33186 4922
rect 33198 4870 33250 4922
rect 33262 4870 33314 4922
rect 33326 4870 33378 4922
rect 3010 4326 3062 4378
rect 3074 4326 3126 4378
rect 3138 4326 3190 4378
rect 3202 4326 3254 4378
rect 3266 4326 3318 4378
rect 33730 4326 33782 4378
rect 33794 4326 33846 4378
rect 33858 4326 33910 4378
rect 33922 4326 33974 4378
rect 33986 4326 34038 4378
rect 2350 3782 2402 3834
rect 2414 3782 2466 3834
rect 2478 3782 2530 3834
rect 2542 3782 2594 3834
rect 2606 3782 2658 3834
rect 33070 3782 33122 3834
rect 33134 3782 33186 3834
rect 33198 3782 33250 3834
rect 33262 3782 33314 3834
rect 33326 3782 33378 3834
rect 3010 3238 3062 3290
rect 3074 3238 3126 3290
rect 3138 3238 3190 3290
rect 3202 3238 3254 3290
rect 3266 3238 3318 3290
rect 33730 3238 33782 3290
rect 33794 3238 33846 3290
rect 33858 3238 33910 3290
rect 33922 3238 33974 3290
rect 33986 3238 34038 3290
rect 2350 2694 2402 2746
rect 2414 2694 2466 2746
rect 2478 2694 2530 2746
rect 2542 2694 2594 2746
rect 2606 2694 2658 2746
rect 33070 2694 33122 2746
rect 33134 2694 33186 2746
rect 33198 2694 33250 2746
rect 33262 2694 33314 2746
rect 33326 2694 33378 2746
rect 3010 2150 3062 2202
rect 3074 2150 3126 2202
rect 3138 2150 3190 2202
rect 3202 2150 3254 2202
rect 3266 2150 3318 2202
rect 33730 2150 33782 2202
rect 33794 2150 33846 2202
rect 33858 2150 33910 2202
rect 33922 2150 33974 2202
rect 33986 2150 34038 2202
<< metal2 >>
rect 938 59200 994 60000
rect 2870 59200 2926 60000
rect 4802 59200 4858 60000
rect 6734 59200 6790 60000
rect 8666 59200 8722 60000
rect 10598 59200 10654 60000
rect 12530 59200 12586 60000
rect 14462 59200 14518 60000
rect 16394 59200 16450 60000
rect 18326 59200 18382 60000
rect 20258 59200 20314 60000
rect 22190 59200 22246 60000
rect 24122 59200 24178 60000
rect 26054 59200 26110 60000
rect 27986 59200 28042 60000
rect 29918 59200 29974 60000
rect 30024 59214 30328 59242
rect 952 57458 980 59200
rect 2884 57526 2912 59200
rect 3010 57692 3318 57701
rect 3010 57690 3016 57692
rect 3072 57690 3096 57692
rect 3152 57690 3176 57692
rect 3232 57690 3256 57692
rect 3312 57690 3318 57692
rect 3072 57638 3074 57690
rect 3254 57638 3256 57690
rect 3010 57636 3016 57638
rect 3072 57636 3096 57638
rect 3152 57636 3176 57638
rect 3232 57636 3256 57638
rect 3312 57636 3318 57638
rect 3010 57627 3318 57636
rect 4816 57526 4844 59200
rect 6748 57594 6776 59200
rect 6736 57588 6788 57594
rect 6736 57530 6788 57536
rect 8680 57526 8708 59200
rect 10612 57526 10640 59200
rect 12544 57526 12572 59200
rect 14476 57526 14504 59200
rect 15292 57588 15344 57594
rect 15292 57530 15344 57536
rect 2872 57520 2924 57526
rect 2872 57462 2924 57468
rect 4804 57520 4856 57526
rect 4804 57462 4856 57468
rect 8668 57520 8720 57526
rect 8668 57462 8720 57468
rect 10600 57520 10652 57526
rect 10600 57462 10652 57468
rect 12532 57520 12584 57526
rect 12532 57462 12584 57468
rect 14464 57520 14516 57526
rect 14464 57462 14516 57468
rect 15200 57520 15252 57526
rect 15200 57462 15252 57468
rect 940 57452 992 57458
rect 940 57394 992 57400
rect 4068 57452 4120 57458
rect 4068 57394 4120 57400
rect 5264 57452 5316 57458
rect 5264 57394 5316 57400
rect 7196 57452 7248 57458
rect 7196 57394 7248 57400
rect 2350 57148 2658 57157
rect 2350 57146 2356 57148
rect 2412 57146 2436 57148
rect 2492 57146 2516 57148
rect 2572 57146 2596 57148
rect 2652 57146 2658 57148
rect 2412 57094 2414 57146
rect 2594 57094 2596 57146
rect 2350 57092 2356 57094
rect 2412 57092 2436 57094
rect 2492 57092 2516 57094
rect 2572 57092 2596 57094
rect 2652 57092 2658 57094
rect 2350 57083 2658 57092
rect 3010 56604 3318 56613
rect 3010 56602 3016 56604
rect 3072 56602 3096 56604
rect 3152 56602 3176 56604
rect 3232 56602 3256 56604
rect 3312 56602 3318 56604
rect 3072 56550 3074 56602
rect 3254 56550 3256 56602
rect 3010 56548 3016 56550
rect 3072 56548 3096 56550
rect 3152 56548 3176 56550
rect 3232 56548 3256 56550
rect 3312 56548 3318 56550
rect 3010 56539 3318 56548
rect 2350 56060 2658 56069
rect 2350 56058 2356 56060
rect 2412 56058 2436 56060
rect 2492 56058 2516 56060
rect 2572 56058 2596 56060
rect 2652 56058 2658 56060
rect 2412 56006 2414 56058
rect 2594 56006 2596 56058
rect 2350 56004 2356 56006
rect 2412 56004 2436 56006
rect 2492 56004 2516 56006
rect 2572 56004 2596 56006
rect 2652 56004 2658 56006
rect 2350 55995 2658 56004
rect 4080 55826 4108 57394
rect 5276 56982 5304 57394
rect 5264 56976 5316 56982
rect 5264 56918 5316 56924
rect 7208 56778 7236 57394
rect 7196 56772 7248 56778
rect 7196 56714 7248 56720
rect 15212 56506 15240 57462
rect 15304 56506 15332 57530
rect 16408 57526 16436 59200
rect 18340 57526 18368 59200
rect 20272 57526 20300 59200
rect 22204 57526 22232 59200
rect 24136 57526 24164 59200
rect 26068 58290 26096 59200
rect 26068 58262 26188 58290
rect 26160 57882 26188 58262
rect 26160 57854 26280 57882
rect 26252 57594 26280 57854
rect 28000 57594 28028 59200
rect 29932 59106 29960 59200
rect 30024 59106 30052 59214
rect 29932 59078 30052 59106
rect 30300 57882 30328 59214
rect 31850 59200 31906 60000
rect 33782 59200 33838 60000
rect 33888 59214 34192 59242
rect 30300 57854 30420 57882
rect 30392 57594 30420 57854
rect 26240 57588 26292 57594
rect 26240 57530 26292 57536
rect 27988 57588 28040 57594
rect 27988 57530 28040 57536
rect 30380 57588 30432 57594
rect 30380 57530 30432 57536
rect 31864 57526 31892 59200
rect 33796 59106 33824 59200
rect 33888 59106 33916 59214
rect 33796 59078 33916 59106
rect 33730 57692 34038 57701
rect 33730 57690 33736 57692
rect 33792 57690 33816 57692
rect 33872 57690 33896 57692
rect 33952 57690 33976 57692
rect 34032 57690 34038 57692
rect 33792 57638 33794 57690
rect 33974 57638 33976 57690
rect 33730 57636 33736 57638
rect 33792 57636 33816 57638
rect 33872 57636 33896 57638
rect 33952 57636 33976 57638
rect 34032 57636 34038 57638
rect 33730 57627 34038 57636
rect 34164 57594 34192 59214
rect 35714 59200 35770 60000
rect 37646 59200 37702 60000
rect 39578 59200 39634 60000
rect 41510 59200 41566 60000
rect 43442 59200 43498 60000
rect 45374 59200 45430 60000
rect 47306 59200 47362 60000
rect 49238 59200 49294 60000
rect 49344 59214 49648 59242
rect 35728 57594 35756 59200
rect 34152 57588 34204 57594
rect 34152 57530 34204 57536
rect 35716 57588 35768 57594
rect 35716 57530 35768 57536
rect 37660 57526 37688 59200
rect 39592 57526 39620 59200
rect 41524 57526 41552 59200
rect 43456 57526 43484 59200
rect 45388 57594 45416 59200
rect 47320 57594 47348 59200
rect 49252 59106 49280 59200
rect 49344 59106 49372 59214
rect 49252 59078 49372 59106
rect 45376 57588 45428 57594
rect 45376 57530 45428 57536
rect 47308 57588 47360 57594
rect 49620 57576 49648 59214
rect 51170 59200 51226 60000
rect 53102 59200 53158 60000
rect 55034 59200 55090 60000
rect 56966 59200 57022 60000
rect 58898 59200 58954 60000
rect 51184 57594 51212 59200
rect 53116 57594 53144 59200
rect 55048 57594 55076 59200
rect 56980 57594 57008 59200
rect 49700 57588 49752 57594
rect 49620 57548 49700 57576
rect 47308 57530 47360 57536
rect 49700 57530 49752 57536
rect 51172 57588 51224 57594
rect 51172 57530 51224 57536
rect 53104 57588 53156 57594
rect 53104 57530 53156 57536
rect 55036 57588 55088 57594
rect 55036 57530 55088 57536
rect 56968 57588 57020 57594
rect 56968 57530 57020 57536
rect 58912 57526 58940 59200
rect 16396 57520 16448 57526
rect 16396 57462 16448 57468
rect 18328 57520 18380 57526
rect 18328 57462 18380 57468
rect 20260 57520 20312 57526
rect 20260 57462 20312 57468
rect 22192 57520 22244 57526
rect 22192 57462 22244 57468
rect 24124 57520 24176 57526
rect 24124 57462 24176 57468
rect 31852 57520 31904 57526
rect 31852 57462 31904 57468
rect 37648 57520 37700 57526
rect 37648 57462 37700 57468
rect 39580 57520 39632 57526
rect 39580 57462 39632 57468
rect 41512 57520 41564 57526
rect 41512 57462 41564 57468
rect 43444 57520 43496 57526
rect 43444 57462 43496 57468
rect 53012 57520 53064 57526
rect 53012 57462 53064 57468
rect 56140 57520 56192 57526
rect 56140 57462 56192 57468
rect 58900 57520 58952 57526
rect 58900 57462 58952 57468
rect 16764 57452 16816 57458
rect 16764 57394 16816 57400
rect 17224 57452 17276 57458
rect 17224 57394 17276 57400
rect 18880 57452 18932 57458
rect 18880 57394 18932 57400
rect 20720 57452 20772 57458
rect 20720 57394 20772 57400
rect 22468 57452 22520 57458
rect 22468 57394 22520 57400
rect 24768 57452 24820 57458
rect 24768 57394 24820 57400
rect 27068 57452 27120 57458
rect 27068 57394 27120 57400
rect 27712 57452 27764 57458
rect 27712 57394 27764 57400
rect 30104 57452 30156 57458
rect 30104 57394 30156 57400
rect 32496 57452 32548 57458
rect 32496 57394 32548 57400
rect 34244 57452 34296 57458
rect 34244 57394 34296 57400
rect 35900 57452 35952 57458
rect 35900 57394 35952 57400
rect 38108 57452 38160 57458
rect 38108 57394 38160 57400
rect 40224 57452 40276 57458
rect 40224 57394 40276 57400
rect 41972 57452 42024 57458
rect 41972 57394 42024 57400
rect 43904 57452 43956 57458
rect 43904 57394 43956 57400
rect 45560 57452 45612 57458
rect 45560 57394 45612 57400
rect 47676 57452 47728 57458
rect 47676 57394 47728 57400
rect 49424 57452 49476 57458
rect 49424 57394 49476 57400
rect 51172 57452 51224 57458
rect 51172 57394 51224 57400
rect 52000 57452 52052 57458
rect 52000 57394 52052 57400
rect 16120 57316 16172 57322
rect 16120 57258 16172 57264
rect 16028 57044 16080 57050
rect 16028 56986 16080 56992
rect 15936 56840 15988 56846
rect 15936 56782 15988 56788
rect 15200 56500 15252 56506
rect 15200 56442 15252 56448
rect 15292 56500 15344 56506
rect 15292 56442 15344 56448
rect 15948 56438 15976 56782
rect 16040 56710 16068 56986
rect 16028 56704 16080 56710
rect 16028 56646 16080 56652
rect 16132 56438 16160 57258
rect 16396 56908 16448 56914
rect 16396 56850 16448 56856
rect 16212 56840 16264 56846
rect 16212 56782 16264 56788
rect 15936 56432 15988 56438
rect 15936 56374 15988 56380
rect 16120 56432 16172 56438
rect 16120 56374 16172 56380
rect 15660 56160 15712 56166
rect 15660 56102 15712 56108
rect 16028 56160 16080 56166
rect 16028 56102 16080 56108
rect 4068 55820 4120 55826
rect 4068 55762 4120 55768
rect 15672 55758 15700 56102
rect 16040 55758 16068 56102
rect 15660 55752 15712 55758
rect 15660 55694 15712 55700
rect 16028 55752 16080 55758
rect 16028 55694 16080 55700
rect 16132 55690 16160 56374
rect 16120 55684 16172 55690
rect 16120 55626 16172 55632
rect 15936 55616 15988 55622
rect 15936 55558 15988 55564
rect 3010 55516 3318 55525
rect 3010 55514 3016 55516
rect 3072 55514 3096 55516
rect 3152 55514 3176 55516
rect 3232 55514 3256 55516
rect 3312 55514 3318 55516
rect 3072 55462 3074 55514
rect 3254 55462 3256 55514
rect 3010 55460 3016 55462
rect 3072 55460 3096 55462
rect 3152 55460 3176 55462
rect 3232 55460 3256 55462
rect 3312 55460 3318 55462
rect 3010 55451 3318 55460
rect 2350 54972 2658 54981
rect 2350 54970 2356 54972
rect 2412 54970 2436 54972
rect 2492 54970 2516 54972
rect 2572 54970 2596 54972
rect 2652 54970 2658 54972
rect 2412 54918 2414 54970
rect 2594 54918 2596 54970
rect 2350 54916 2356 54918
rect 2412 54916 2436 54918
rect 2492 54916 2516 54918
rect 2572 54916 2596 54918
rect 2652 54916 2658 54918
rect 2350 54907 2658 54916
rect 15948 54534 15976 55558
rect 15936 54528 15988 54534
rect 15936 54470 15988 54476
rect 3010 54428 3318 54437
rect 3010 54426 3016 54428
rect 3072 54426 3096 54428
rect 3152 54426 3176 54428
rect 3232 54426 3256 54428
rect 3312 54426 3318 54428
rect 3072 54374 3074 54426
rect 3254 54374 3256 54426
rect 3010 54372 3016 54374
rect 3072 54372 3096 54374
rect 3152 54372 3176 54374
rect 3232 54372 3256 54374
rect 3312 54372 3318 54374
rect 3010 54363 3318 54372
rect 16224 53990 16252 56782
rect 16408 56302 16436 56850
rect 16672 56840 16724 56846
rect 16672 56782 16724 56788
rect 16396 56296 16448 56302
rect 16396 56238 16448 56244
rect 16684 55962 16712 56782
rect 16776 56506 16804 57394
rect 16856 57384 16908 57390
rect 16856 57326 16908 57332
rect 16868 56846 16896 57326
rect 17132 56908 17184 56914
rect 17132 56850 17184 56856
rect 16856 56840 16908 56846
rect 16856 56782 16908 56788
rect 16764 56500 16816 56506
rect 16764 56442 16816 56448
rect 16868 56438 16896 56782
rect 17144 56710 17172 56850
rect 16948 56704 17000 56710
rect 16948 56646 17000 56652
rect 17132 56704 17184 56710
rect 17132 56646 17184 56652
rect 16856 56432 16908 56438
rect 16856 56374 16908 56380
rect 16672 55956 16724 55962
rect 16672 55898 16724 55904
rect 16764 55616 16816 55622
rect 16764 55558 16816 55564
rect 16776 55282 16804 55558
rect 16868 55350 16896 56374
rect 16960 55758 16988 56646
rect 16948 55752 17000 55758
rect 16948 55694 17000 55700
rect 16948 55616 17000 55622
rect 17144 55570 17172 56646
rect 17236 56370 17264 57394
rect 17316 56908 17368 56914
rect 17316 56850 17368 56856
rect 17868 56908 17920 56914
rect 17868 56850 17920 56856
rect 17224 56364 17276 56370
rect 17224 56306 17276 56312
rect 17328 56302 17356 56850
rect 17408 56704 17460 56710
rect 17408 56646 17460 56652
rect 17420 56545 17448 56646
rect 17406 56536 17462 56545
rect 17406 56471 17462 56480
rect 17776 56500 17828 56506
rect 17776 56442 17828 56448
rect 17316 56296 17368 56302
rect 17316 56238 17368 56244
rect 17328 55826 17356 56238
rect 17592 56228 17644 56234
rect 17592 56170 17644 56176
rect 17500 56160 17552 56166
rect 17500 56102 17552 56108
rect 17316 55820 17368 55826
rect 17316 55762 17368 55768
rect 17224 55752 17276 55758
rect 17224 55694 17276 55700
rect 17236 55622 17264 55694
rect 17224 55616 17276 55622
rect 17000 55564 17172 55570
rect 16948 55558 17172 55564
rect 16960 55542 17172 55558
rect 17222 55584 17224 55593
rect 17276 55584 17278 55593
rect 17222 55519 17278 55528
rect 16856 55344 16908 55350
rect 17328 55321 17356 55762
rect 16856 55286 16908 55292
rect 16946 55312 17002 55321
rect 16764 55276 16816 55282
rect 16946 55247 17002 55256
rect 17314 55312 17370 55321
rect 17512 55282 17540 56102
rect 17604 55826 17632 56170
rect 17592 55820 17644 55826
rect 17592 55762 17644 55768
rect 17788 55758 17816 56442
rect 17880 55894 17908 56850
rect 18144 56840 18196 56846
rect 18144 56782 18196 56788
rect 17960 56772 18012 56778
rect 17960 56714 18012 56720
rect 17868 55888 17920 55894
rect 17868 55830 17920 55836
rect 17776 55752 17828 55758
rect 17776 55694 17828 55700
rect 17314 55247 17370 55256
rect 17500 55276 17552 55282
rect 16764 55218 16816 55224
rect 16960 55214 16988 55247
rect 17500 55218 17552 55224
rect 16948 55208 17000 55214
rect 16948 55150 17000 55156
rect 16212 53984 16264 53990
rect 16212 53926 16264 53932
rect 2350 53884 2658 53893
rect 2350 53882 2356 53884
rect 2412 53882 2436 53884
rect 2492 53882 2516 53884
rect 2572 53882 2596 53884
rect 2652 53882 2658 53884
rect 2412 53830 2414 53882
rect 2594 53830 2596 53882
rect 2350 53828 2356 53830
rect 2412 53828 2436 53830
rect 2492 53828 2516 53830
rect 2572 53828 2596 53830
rect 2652 53828 2658 53830
rect 2350 53819 2658 53828
rect 17788 53786 17816 55694
rect 17972 55214 18000 56714
rect 18156 55962 18184 56782
rect 18604 56704 18656 56710
rect 18604 56646 18656 56652
rect 18328 56160 18380 56166
rect 18328 56102 18380 56108
rect 18144 55956 18196 55962
rect 18144 55898 18196 55904
rect 18340 55758 18368 56102
rect 18616 55826 18644 56646
rect 18892 56370 18920 57394
rect 19524 56840 19576 56846
rect 19524 56782 19576 56788
rect 19248 56500 19300 56506
rect 19300 56460 19380 56488
rect 19248 56442 19300 56448
rect 18880 56364 18932 56370
rect 18880 56306 18932 56312
rect 18696 56296 18748 56302
rect 18696 56238 18748 56244
rect 18708 55962 18736 56238
rect 18892 56234 18920 56306
rect 18880 56228 18932 56234
rect 18880 56170 18932 56176
rect 19352 56166 19380 56460
rect 19432 56364 19484 56370
rect 19432 56306 19484 56312
rect 19444 56234 19472 56306
rect 19432 56228 19484 56234
rect 19432 56170 19484 56176
rect 19340 56160 19392 56166
rect 19340 56102 19392 56108
rect 18696 55956 18748 55962
rect 18696 55898 18748 55904
rect 19340 55888 19392 55894
rect 19340 55830 19392 55836
rect 18604 55820 18656 55826
rect 18604 55762 18656 55768
rect 18328 55752 18380 55758
rect 18328 55694 18380 55700
rect 17960 55208 18012 55214
rect 17960 55150 18012 55156
rect 19352 54806 19380 55830
rect 19340 54800 19392 54806
rect 19340 54742 19392 54748
rect 17776 53780 17828 53786
rect 17776 53722 17828 53728
rect 3010 53340 3318 53349
rect 3010 53338 3016 53340
rect 3072 53338 3096 53340
rect 3152 53338 3176 53340
rect 3232 53338 3256 53340
rect 3312 53338 3318 53340
rect 3072 53286 3074 53338
rect 3254 53286 3256 53338
rect 3010 53284 3016 53286
rect 3072 53284 3096 53286
rect 3152 53284 3176 53286
rect 3232 53284 3256 53286
rect 3312 53284 3318 53286
rect 3010 53275 3318 53284
rect 19444 53242 19472 56170
rect 19536 55826 19564 56782
rect 19890 56536 19946 56545
rect 19890 56471 19946 56480
rect 19904 56166 19932 56471
rect 19984 56296 20036 56302
rect 19984 56238 20036 56244
rect 19616 56160 19668 56166
rect 19616 56102 19668 56108
rect 19708 56160 19760 56166
rect 19708 56102 19760 56108
rect 19892 56160 19944 56166
rect 19892 56102 19944 56108
rect 19628 55894 19656 56102
rect 19616 55888 19668 55894
rect 19616 55830 19668 55836
rect 19524 55820 19576 55826
rect 19524 55762 19576 55768
rect 19720 55758 19748 56102
rect 19800 55956 19852 55962
rect 19800 55898 19852 55904
rect 19708 55752 19760 55758
rect 19708 55694 19760 55700
rect 19616 55684 19668 55690
rect 19616 55626 19668 55632
rect 19628 55593 19656 55626
rect 19614 55584 19670 55593
rect 19614 55519 19670 55528
rect 19812 55418 19840 55898
rect 19708 55412 19760 55418
rect 19708 55354 19760 55360
rect 19800 55412 19852 55418
rect 19800 55354 19852 55360
rect 19616 55344 19668 55350
rect 19616 55286 19668 55292
rect 19628 54330 19656 55286
rect 19720 55214 19748 55354
rect 19720 55208 19944 55214
rect 19720 55186 19892 55208
rect 19892 55150 19944 55156
rect 19996 55078 20024 56238
rect 20732 56166 20760 57394
rect 21272 57044 21324 57050
rect 21272 56986 21324 56992
rect 20812 56976 20864 56982
rect 20812 56918 20864 56924
rect 20720 56160 20772 56166
rect 20720 56102 20772 56108
rect 20444 55888 20496 55894
rect 20444 55830 20496 55836
rect 20534 55856 20590 55865
rect 19984 55072 20036 55078
rect 19984 55014 20036 55020
rect 20456 54874 20484 55830
rect 20534 55791 20536 55800
rect 20588 55791 20590 55800
rect 20536 55762 20588 55768
rect 20628 55616 20680 55622
rect 20628 55558 20680 55564
rect 20444 54868 20496 54874
rect 20444 54810 20496 54816
rect 19616 54324 19668 54330
rect 19616 54266 19668 54272
rect 19432 53236 19484 53242
rect 19432 53178 19484 53184
rect 20640 53038 20668 55558
rect 20824 54126 20852 56918
rect 20904 56772 20956 56778
rect 20904 56714 20956 56720
rect 20916 56438 20944 56714
rect 21284 56438 21312 56986
rect 22480 56846 22508 57394
rect 22192 56840 22244 56846
rect 22192 56782 22244 56788
rect 22468 56840 22520 56846
rect 22468 56782 22520 56788
rect 20904 56432 20956 56438
rect 20904 56374 20956 56380
rect 21272 56432 21324 56438
rect 21272 56374 21324 56380
rect 20916 55350 20944 56374
rect 21824 56160 21876 56166
rect 21824 56102 21876 56108
rect 22100 56160 22152 56166
rect 22204 56148 22232 56782
rect 22480 56370 22508 56782
rect 22560 56704 22612 56710
rect 22560 56646 22612 56652
rect 23664 56704 23716 56710
rect 23664 56646 23716 56652
rect 22468 56364 22520 56370
rect 22468 56306 22520 56312
rect 22284 56296 22336 56302
rect 22284 56238 22336 56244
rect 22152 56120 22232 56148
rect 22100 56102 22152 56108
rect 20904 55344 20956 55350
rect 20904 55286 20956 55292
rect 21836 55214 21864 56102
rect 21916 55888 21968 55894
rect 21914 55856 21916 55865
rect 21968 55856 21970 55865
rect 22112 55826 22140 56102
rect 21914 55791 21970 55800
rect 22100 55820 22152 55826
rect 22100 55762 22152 55768
rect 22008 55752 22060 55758
rect 22008 55694 22060 55700
rect 22020 55350 22048 55694
rect 22112 55418 22140 55762
rect 22100 55412 22152 55418
rect 22100 55354 22152 55360
rect 22008 55344 22060 55350
rect 22008 55286 22060 55292
rect 21824 55208 21876 55214
rect 21824 55150 21876 55156
rect 22020 54602 22048 55286
rect 22112 55282 22140 55354
rect 22296 55282 22324 56238
rect 22376 56160 22428 56166
rect 22376 56102 22428 56108
rect 22388 55962 22416 56102
rect 22376 55956 22428 55962
rect 22376 55898 22428 55904
rect 22480 55842 22508 56306
rect 22388 55814 22508 55842
rect 22388 55622 22416 55814
rect 22376 55616 22428 55622
rect 22376 55558 22428 55564
rect 22468 55412 22520 55418
rect 22468 55354 22520 55360
rect 22100 55276 22152 55282
rect 22100 55218 22152 55224
rect 22284 55276 22336 55282
rect 22284 55218 22336 55224
rect 22480 54738 22508 55354
rect 22468 54732 22520 54738
rect 22468 54674 22520 54680
rect 22008 54596 22060 54602
rect 22008 54538 22060 54544
rect 22020 54262 22048 54538
rect 21088 54256 21140 54262
rect 21088 54198 21140 54204
rect 22008 54256 22060 54262
rect 22008 54198 22060 54204
rect 20812 54120 20864 54126
rect 20812 54062 20864 54068
rect 21100 53582 21128 54198
rect 22480 54126 22508 54674
rect 22468 54120 22520 54126
rect 22468 54062 22520 54068
rect 22480 53650 22508 54062
rect 22468 53644 22520 53650
rect 22468 53586 22520 53592
rect 21088 53576 21140 53582
rect 21088 53518 21140 53524
rect 21100 53174 21128 53518
rect 21088 53168 21140 53174
rect 21088 53110 21140 53116
rect 22480 53106 22508 53586
rect 22572 53514 22600 56646
rect 23676 56506 23704 56646
rect 24780 56506 24808 57394
rect 27080 56846 27108 57394
rect 27068 56840 27120 56846
rect 27068 56782 27120 56788
rect 26516 56704 26568 56710
rect 26516 56646 26568 56652
rect 26528 56506 26556 56646
rect 23664 56500 23716 56506
rect 23664 56442 23716 56448
rect 24768 56500 24820 56506
rect 24768 56442 24820 56448
rect 26516 56500 26568 56506
rect 26516 56442 26568 56448
rect 23756 56432 23808 56438
rect 23756 56374 23808 56380
rect 22744 56160 22796 56166
rect 22744 56102 22796 56108
rect 22756 55690 22784 56102
rect 23768 55894 23796 56374
rect 24780 55978 24808 56442
rect 27080 56438 27108 56782
rect 27160 56704 27212 56710
rect 27160 56646 27212 56652
rect 27068 56432 27120 56438
rect 27068 56374 27120 56380
rect 25044 56160 25096 56166
rect 25044 56102 25096 56108
rect 26976 56160 27028 56166
rect 26976 56102 27028 56108
rect 24688 55950 24808 55978
rect 24688 55894 24716 55950
rect 23756 55888 23808 55894
rect 23756 55830 23808 55836
rect 24676 55888 24728 55894
rect 24676 55830 24728 55836
rect 24768 55820 24820 55826
rect 24768 55762 24820 55768
rect 23848 55752 23900 55758
rect 23848 55694 23900 55700
rect 22744 55684 22796 55690
rect 22744 55626 22796 55632
rect 23020 55616 23072 55622
rect 22834 55584 22890 55593
rect 23020 55558 23072 55564
rect 23112 55616 23164 55622
rect 23112 55558 23164 55564
rect 22834 55519 22890 55528
rect 22848 55282 22876 55519
rect 23032 55282 23060 55558
rect 23124 55350 23152 55558
rect 23112 55344 23164 55350
rect 23112 55286 23164 55292
rect 22836 55276 22888 55282
rect 22836 55218 22888 55224
rect 23020 55276 23072 55282
rect 23020 55218 23072 55224
rect 23296 55072 23348 55078
rect 23296 55014 23348 55020
rect 23308 54874 23336 55014
rect 23296 54868 23348 54874
rect 23296 54810 23348 54816
rect 23860 54670 23888 55694
rect 24492 55616 24544 55622
rect 24492 55558 24544 55564
rect 24504 55350 24532 55558
rect 24492 55344 24544 55350
rect 24492 55286 24544 55292
rect 24780 55214 24808 55762
rect 25056 55350 25084 56102
rect 26988 55826 27016 56102
rect 26976 55820 27028 55826
rect 26976 55762 27028 55768
rect 26240 55752 26292 55758
rect 26240 55694 26292 55700
rect 26252 55400 26280 55694
rect 26424 55684 26476 55690
rect 26424 55626 26476 55632
rect 26332 55412 26384 55418
rect 26252 55372 26332 55400
rect 25044 55344 25096 55350
rect 25044 55286 25096 55292
rect 24768 55208 24820 55214
rect 24768 55150 24820 55156
rect 26252 54806 26280 55372
rect 26332 55354 26384 55360
rect 26436 55350 26464 55626
rect 27080 55418 27108 56374
rect 27172 56370 27200 56646
rect 27724 56438 27752 57394
rect 27804 56840 27856 56846
rect 27804 56782 27856 56788
rect 28172 56840 28224 56846
rect 28172 56782 28224 56788
rect 27816 56506 27844 56782
rect 27896 56704 27948 56710
rect 27896 56646 27948 56652
rect 27804 56500 27856 56506
rect 27804 56442 27856 56448
rect 27712 56432 27764 56438
rect 27712 56374 27764 56380
rect 27160 56364 27212 56370
rect 27160 56306 27212 56312
rect 27724 55894 27752 56374
rect 27712 55888 27764 55894
rect 27712 55830 27764 55836
rect 27804 55684 27856 55690
rect 27804 55626 27856 55632
rect 27068 55412 27120 55418
rect 27068 55354 27120 55360
rect 27816 55350 27844 55626
rect 26424 55344 26476 55350
rect 26424 55286 26476 55292
rect 27804 55344 27856 55350
rect 27804 55286 27856 55292
rect 26516 55276 26568 55282
rect 26516 55218 26568 55224
rect 26240 54800 26292 54806
rect 26240 54742 26292 54748
rect 23848 54664 23900 54670
rect 23848 54606 23900 54612
rect 26528 53786 26556 55218
rect 27908 54738 27936 56646
rect 28184 56506 28212 56782
rect 28172 56500 28224 56506
rect 28172 56442 28224 56448
rect 30116 56438 30144 57394
rect 32508 56506 32536 57394
rect 33070 57148 33378 57157
rect 33070 57146 33076 57148
rect 33132 57146 33156 57148
rect 33212 57146 33236 57148
rect 33292 57146 33316 57148
rect 33372 57146 33378 57148
rect 33132 57094 33134 57146
rect 33314 57094 33316 57146
rect 33070 57092 33076 57094
rect 33132 57092 33156 57094
rect 33212 57092 33236 57094
rect 33292 57092 33316 57094
rect 33372 57092 33378 57094
rect 33070 57083 33378 57092
rect 33730 56604 34038 56613
rect 33730 56602 33736 56604
rect 33792 56602 33816 56604
rect 33872 56602 33896 56604
rect 33952 56602 33976 56604
rect 34032 56602 34038 56604
rect 33792 56550 33794 56602
rect 33974 56550 33976 56602
rect 33730 56548 33736 56550
rect 33792 56548 33816 56550
rect 33872 56548 33896 56550
rect 33952 56548 33976 56550
rect 34032 56548 34038 56550
rect 33730 56539 34038 56548
rect 32220 56500 32272 56506
rect 32220 56442 32272 56448
rect 32496 56500 32548 56506
rect 32496 56442 32548 56448
rect 30104 56432 30156 56438
rect 30104 56374 30156 56380
rect 28724 56296 28776 56302
rect 28724 56238 28776 56244
rect 28080 56160 28132 56166
rect 28080 56102 28132 56108
rect 28092 55758 28120 56102
rect 28736 55894 28764 56238
rect 28724 55888 28776 55894
rect 28724 55830 28776 55836
rect 30116 55826 30144 56374
rect 32232 56302 32260 56442
rect 34256 56302 34284 57394
rect 35912 56506 35940 57394
rect 38120 56506 38148 57394
rect 40236 56506 40264 57394
rect 35900 56500 35952 56506
rect 35900 56442 35952 56448
rect 38108 56500 38160 56506
rect 38108 56442 38160 56448
rect 40224 56500 40276 56506
rect 40224 56442 40276 56448
rect 32220 56296 32272 56302
rect 32220 56238 32272 56244
rect 32680 56296 32732 56302
rect 32680 56238 32732 56244
rect 34244 56296 34296 56302
rect 34244 56238 34296 56244
rect 30104 55820 30156 55826
rect 30104 55762 30156 55768
rect 28080 55752 28132 55758
rect 28080 55694 28132 55700
rect 28448 55616 28500 55622
rect 28448 55558 28500 55564
rect 29552 55616 29604 55622
rect 29552 55558 29604 55564
rect 28460 55350 28488 55558
rect 28448 55344 28500 55350
rect 28448 55286 28500 55292
rect 29564 55282 29592 55558
rect 29552 55276 29604 55282
rect 29552 55218 29604 55224
rect 27896 54732 27948 54738
rect 27896 54674 27948 54680
rect 29564 54670 29592 55218
rect 30116 54874 30144 55762
rect 32036 55412 32088 55418
rect 32232 55400 32260 56238
rect 32404 56160 32456 56166
rect 32404 56102 32456 56108
rect 32088 55372 32260 55400
rect 32036 55354 32088 55360
rect 32416 55350 32444 56102
rect 32692 55894 32720 56238
rect 33070 56060 33378 56069
rect 33070 56058 33076 56060
rect 33132 56058 33156 56060
rect 33212 56058 33236 56060
rect 33292 56058 33316 56060
rect 33372 56058 33378 56060
rect 33132 56006 33134 56058
rect 33314 56006 33316 56058
rect 33070 56004 33076 56006
rect 33132 56004 33156 56006
rect 33212 56004 33236 56006
rect 33292 56004 33316 56006
rect 33372 56004 33378 56006
rect 33070 55995 33378 56004
rect 32680 55888 32732 55894
rect 32680 55830 32732 55836
rect 33416 55616 33468 55622
rect 33416 55558 33468 55564
rect 33428 55350 33456 55558
rect 33730 55516 34038 55525
rect 33730 55514 33736 55516
rect 33792 55514 33816 55516
rect 33872 55514 33896 55516
rect 33952 55514 33976 55516
rect 34032 55514 34038 55516
rect 33792 55462 33794 55514
rect 33974 55462 33976 55514
rect 33730 55460 33736 55462
rect 33792 55460 33816 55462
rect 33872 55460 33896 55462
rect 33952 55460 33976 55462
rect 34032 55460 34038 55462
rect 33730 55451 34038 55460
rect 32404 55344 32456 55350
rect 32404 55286 32456 55292
rect 33416 55344 33468 55350
rect 33416 55286 33468 55292
rect 34256 55078 34284 56238
rect 34796 56160 34848 56166
rect 34796 56102 34848 56108
rect 34808 55214 34836 56102
rect 35532 55616 35584 55622
rect 35532 55558 35584 55564
rect 35544 55350 35572 55558
rect 35912 55418 35940 56442
rect 36268 56364 36320 56370
rect 36268 56306 36320 56312
rect 36176 55684 36228 55690
rect 36176 55626 36228 55632
rect 35900 55412 35952 55418
rect 35900 55354 35952 55360
rect 35532 55344 35584 55350
rect 35532 55286 35584 55292
rect 34796 55208 34848 55214
rect 34796 55150 34848 55156
rect 34244 55072 34296 55078
rect 34244 55014 34296 55020
rect 33070 54972 33378 54981
rect 33070 54970 33076 54972
rect 33132 54970 33156 54972
rect 33212 54970 33236 54972
rect 33292 54970 33316 54972
rect 33372 54970 33378 54972
rect 33132 54918 33134 54970
rect 33314 54918 33316 54970
rect 33070 54916 33076 54918
rect 33132 54916 33156 54918
rect 33212 54916 33236 54918
rect 33292 54916 33316 54918
rect 33372 54916 33378 54918
rect 33070 54907 33378 54916
rect 30104 54868 30156 54874
rect 30104 54810 30156 54816
rect 29552 54664 29604 54670
rect 29552 54606 29604 54612
rect 36188 54602 36216 55626
rect 36280 54874 36308 56306
rect 37740 56160 37792 56166
rect 37740 56102 37792 56108
rect 38660 56160 38712 56166
rect 38660 56102 38712 56108
rect 40132 56160 40184 56166
rect 40132 56102 40184 56108
rect 37280 55344 37332 55350
rect 37280 55286 37332 55292
rect 36268 54868 36320 54874
rect 36268 54810 36320 54816
rect 37292 54602 37320 55286
rect 37752 54738 37780 56102
rect 38016 55684 38068 55690
rect 38016 55626 38068 55632
rect 37924 55412 37976 55418
rect 37924 55354 37976 55360
rect 37936 55282 37964 55354
rect 37924 55276 37976 55282
rect 37924 55218 37976 55224
rect 38028 55214 38056 55626
rect 38476 55412 38528 55418
rect 38476 55354 38528 55360
rect 38488 55214 38516 55354
rect 38672 55298 38700 56102
rect 38028 55186 38148 55214
rect 38016 55072 38068 55078
rect 38016 55014 38068 55020
rect 38028 54738 38056 55014
rect 37740 54732 37792 54738
rect 37740 54674 37792 54680
rect 38016 54732 38068 54738
rect 38016 54674 38068 54680
rect 36176 54596 36228 54602
rect 36176 54538 36228 54544
rect 37280 54596 37332 54602
rect 37280 54538 37332 54544
rect 27804 54528 27856 54534
rect 27804 54470 27856 54476
rect 26516 53780 26568 53786
rect 26516 53722 26568 53728
rect 27816 53582 27844 54470
rect 33730 54428 34038 54437
rect 33730 54426 33736 54428
rect 33792 54426 33816 54428
rect 33872 54426 33896 54428
rect 33952 54426 33976 54428
rect 34032 54426 34038 54428
rect 33792 54374 33794 54426
rect 33974 54374 33976 54426
rect 33730 54372 33736 54374
rect 33792 54372 33816 54374
rect 33872 54372 33896 54374
rect 33952 54372 33976 54374
rect 34032 54372 34038 54374
rect 33730 54363 34038 54372
rect 33070 53884 33378 53893
rect 33070 53882 33076 53884
rect 33132 53882 33156 53884
rect 33212 53882 33236 53884
rect 33292 53882 33316 53884
rect 33372 53882 33378 53884
rect 33132 53830 33134 53882
rect 33314 53830 33316 53882
rect 33070 53828 33076 53830
rect 33132 53828 33156 53830
rect 33212 53828 33236 53830
rect 33292 53828 33316 53830
rect 33372 53828 33378 53830
rect 33070 53819 33378 53828
rect 27804 53576 27856 53582
rect 27804 53518 27856 53524
rect 22560 53508 22612 53514
rect 22560 53450 22612 53456
rect 33730 53340 34038 53349
rect 33730 53338 33736 53340
rect 33792 53338 33816 53340
rect 33872 53338 33896 53340
rect 33952 53338 33976 53340
rect 34032 53338 34038 53340
rect 33792 53286 33794 53338
rect 33974 53286 33976 53338
rect 33730 53284 33736 53286
rect 33792 53284 33816 53286
rect 33872 53284 33896 53286
rect 33952 53284 33976 53286
rect 34032 53284 34038 53286
rect 33730 53275 34038 53284
rect 22468 53100 22520 53106
rect 22468 53042 22520 53048
rect 20628 53032 20680 53038
rect 20628 52974 20680 52980
rect 2350 52796 2658 52805
rect 2350 52794 2356 52796
rect 2412 52794 2436 52796
rect 2492 52794 2516 52796
rect 2572 52794 2596 52796
rect 2652 52794 2658 52796
rect 2412 52742 2414 52794
rect 2594 52742 2596 52794
rect 2350 52740 2356 52742
rect 2412 52740 2436 52742
rect 2492 52740 2516 52742
rect 2572 52740 2596 52742
rect 2652 52740 2658 52742
rect 2350 52731 2658 52740
rect 33070 52796 33378 52805
rect 33070 52794 33076 52796
rect 33132 52794 33156 52796
rect 33212 52794 33236 52796
rect 33292 52794 33316 52796
rect 33372 52794 33378 52796
rect 33132 52742 33134 52794
rect 33314 52742 33316 52794
rect 33070 52740 33076 52742
rect 33132 52740 33156 52742
rect 33212 52740 33236 52742
rect 33292 52740 33316 52742
rect 33372 52740 33378 52742
rect 33070 52731 33378 52740
rect 3010 52252 3318 52261
rect 3010 52250 3016 52252
rect 3072 52250 3096 52252
rect 3152 52250 3176 52252
rect 3232 52250 3256 52252
rect 3312 52250 3318 52252
rect 3072 52198 3074 52250
rect 3254 52198 3256 52250
rect 3010 52196 3016 52198
rect 3072 52196 3096 52198
rect 3152 52196 3176 52198
rect 3232 52196 3256 52198
rect 3312 52196 3318 52198
rect 3010 52187 3318 52196
rect 33730 52252 34038 52261
rect 33730 52250 33736 52252
rect 33792 52250 33816 52252
rect 33872 52250 33896 52252
rect 33952 52250 33976 52252
rect 34032 52250 34038 52252
rect 33792 52198 33794 52250
rect 33974 52198 33976 52250
rect 33730 52196 33736 52198
rect 33792 52196 33816 52198
rect 33872 52196 33896 52198
rect 33952 52196 33976 52198
rect 34032 52196 34038 52198
rect 33730 52187 34038 52196
rect 2350 51708 2658 51717
rect 2350 51706 2356 51708
rect 2412 51706 2436 51708
rect 2492 51706 2516 51708
rect 2572 51706 2596 51708
rect 2652 51706 2658 51708
rect 2412 51654 2414 51706
rect 2594 51654 2596 51706
rect 2350 51652 2356 51654
rect 2412 51652 2436 51654
rect 2492 51652 2516 51654
rect 2572 51652 2596 51654
rect 2652 51652 2658 51654
rect 2350 51643 2658 51652
rect 33070 51708 33378 51717
rect 33070 51706 33076 51708
rect 33132 51706 33156 51708
rect 33212 51706 33236 51708
rect 33292 51706 33316 51708
rect 33372 51706 33378 51708
rect 33132 51654 33134 51706
rect 33314 51654 33316 51706
rect 33070 51652 33076 51654
rect 33132 51652 33156 51654
rect 33212 51652 33236 51654
rect 33292 51652 33316 51654
rect 33372 51652 33378 51654
rect 33070 51643 33378 51652
rect 3010 51164 3318 51173
rect 3010 51162 3016 51164
rect 3072 51162 3096 51164
rect 3152 51162 3176 51164
rect 3232 51162 3256 51164
rect 3312 51162 3318 51164
rect 3072 51110 3074 51162
rect 3254 51110 3256 51162
rect 3010 51108 3016 51110
rect 3072 51108 3096 51110
rect 3152 51108 3176 51110
rect 3232 51108 3256 51110
rect 3312 51108 3318 51110
rect 3010 51099 3318 51108
rect 33730 51164 34038 51173
rect 33730 51162 33736 51164
rect 33792 51162 33816 51164
rect 33872 51162 33896 51164
rect 33952 51162 33976 51164
rect 34032 51162 34038 51164
rect 33792 51110 33794 51162
rect 33974 51110 33976 51162
rect 33730 51108 33736 51110
rect 33792 51108 33816 51110
rect 33872 51108 33896 51110
rect 33952 51108 33976 51110
rect 34032 51108 34038 51110
rect 33730 51099 34038 51108
rect 2350 50620 2658 50629
rect 2350 50618 2356 50620
rect 2412 50618 2436 50620
rect 2492 50618 2516 50620
rect 2572 50618 2596 50620
rect 2652 50618 2658 50620
rect 2412 50566 2414 50618
rect 2594 50566 2596 50618
rect 2350 50564 2356 50566
rect 2412 50564 2436 50566
rect 2492 50564 2516 50566
rect 2572 50564 2596 50566
rect 2652 50564 2658 50566
rect 2350 50555 2658 50564
rect 33070 50620 33378 50629
rect 33070 50618 33076 50620
rect 33132 50618 33156 50620
rect 33212 50618 33236 50620
rect 33292 50618 33316 50620
rect 33372 50618 33378 50620
rect 33132 50566 33134 50618
rect 33314 50566 33316 50618
rect 33070 50564 33076 50566
rect 33132 50564 33156 50566
rect 33212 50564 33236 50566
rect 33292 50564 33316 50566
rect 33372 50564 33378 50566
rect 33070 50555 33378 50564
rect 3010 50076 3318 50085
rect 3010 50074 3016 50076
rect 3072 50074 3096 50076
rect 3152 50074 3176 50076
rect 3232 50074 3256 50076
rect 3312 50074 3318 50076
rect 3072 50022 3074 50074
rect 3254 50022 3256 50074
rect 3010 50020 3016 50022
rect 3072 50020 3096 50022
rect 3152 50020 3176 50022
rect 3232 50020 3256 50022
rect 3312 50020 3318 50022
rect 3010 50011 3318 50020
rect 33730 50076 34038 50085
rect 33730 50074 33736 50076
rect 33792 50074 33816 50076
rect 33872 50074 33896 50076
rect 33952 50074 33976 50076
rect 34032 50074 34038 50076
rect 33792 50022 33794 50074
rect 33974 50022 33976 50074
rect 33730 50020 33736 50022
rect 33792 50020 33816 50022
rect 33872 50020 33896 50022
rect 33952 50020 33976 50022
rect 34032 50020 34038 50022
rect 33730 50011 34038 50020
rect 2350 49532 2658 49541
rect 2350 49530 2356 49532
rect 2412 49530 2436 49532
rect 2492 49530 2516 49532
rect 2572 49530 2596 49532
rect 2652 49530 2658 49532
rect 2412 49478 2414 49530
rect 2594 49478 2596 49530
rect 2350 49476 2356 49478
rect 2412 49476 2436 49478
rect 2492 49476 2516 49478
rect 2572 49476 2596 49478
rect 2652 49476 2658 49478
rect 2350 49467 2658 49476
rect 33070 49532 33378 49541
rect 33070 49530 33076 49532
rect 33132 49530 33156 49532
rect 33212 49530 33236 49532
rect 33292 49530 33316 49532
rect 33372 49530 33378 49532
rect 33132 49478 33134 49530
rect 33314 49478 33316 49530
rect 33070 49476 33076 49478
rect 33132 49476 33156 49478
rect 33212 49476 33236 49478
rect 33292 49476 33316 49478
rect 33372 49476 33378 49478
rect 33070 49467 33378 49476
rect 3010 48988 3318 48997
rect 3010 48986 3016 48988
rect 3072 48986 3096 48988
rect 3152 48986 3176 48988
rect 3232 48986 3256 48988
rect 3312 48986 3318 48988
rect 3072 48934 3074 48986
rect 3254 48934 3256 48986
rect 3010 48932 3016 48934
rect 3072 48932 3096 48934
rect 3152 48932 3176 48934
rect 3232 48932 3256 48934
rect 3312 48932 3318 48934
rect 3010 48923 3318 48932
rect 33730 48988 34038 48997
rect 33730 48986 33736 48988
rect 33792 48986 33816 48988
rect 33872 48986 33896 48988
rect 33952 48986 33976 48988
rect 34032 48986 34038 48988
rect 33792 48934 33794 48986
rect 33974 48934 33976 48986
rect 33730 48932 33736 48934
rect 33792 48932 33816 48934
rect 33872 48932 33896 48934
rect 33952 48932 33976 48934
rect 34032 48932 34038 48934
rect 33730 48923 34038 48932
rect 2350 48444 2658 48453
rect 2350 48442 2356 48444
rect 2412 48442 2436 48444
rect 2492 48442 2516 48444
rect 2572 48442 2596 48444
rect 2652 48442 2658 48444
rect 2412 48390 2414 48442
rect 2594 48390 2596 48442
rect 2350 48388 2356 48390
rect 2412 48388 2436 48390
rect 2492 48388 2516 48390
rect 2572 48388 2596 48390
rect 2652 48388 2658 48390
rect 2350 48379 2658 48388
rect 33070 48444 33378 48453
rect 33070 48442 33076 48444
rect 33132 48442 33156 48444
rect 33212 48442 33236 48444
rect 33292 48442 33316 48444
rect 33372 48442 33378 48444
rect 33132 48390 33134 48442
rect 33314 48390 33316 48442
rect 33070 48388 33076 48390
rect 33132 48388 33156 48390
rect 33212 48388 33236 48390
rect 33292 48388 33316 48390
rect 33372 48388 33378 48390
rect 33070 48379 33378 48388
rect 3010 47900 3318 47909
rect 3010 47898 3016 47900
rect 3072 47898 3096 47900
rect 3152 47898 3176 47900
rect 3232 47898 3256 47900
rect 3312 47898 3318 47900
rect 3072 47846 3074 47898
rect 3254 47846 3256 47898
rect 3010 47844 3016 47846
rect 3072 47844 3096 47846
rect 3152 47844 3176 47846
rect 3232 47844 3256 47846
rect 3312 47844 3318 47846
rect 3010 47835 3318 47844
rect 33730 47900 34038 47909
rect 33730 47898 33736 47900
rect 33792 47898 33816 47900
rect 33872 47898 33896 47900
rect 33952 47898 33976 47900
rect 34032 47898 34038 47900
rect 33792 47846 33794 47898
rect 33974 47846 33976 47898
rect 33730 47844 33736 47846
rect 33792 47844 33816 47846
rect 33872 47844 33896 47846
rect 33952 47844 33976 47846
rect 34032 47844 34038 47846
rect 33730 47835 34038 47844
rect 2350 47356 2658 47365
rect 2350 47354 2356 47356
rect 2412 47354 2436 47356
rect 2492 47354 2516 47356
rect 2572 47354 2596 47356
rect 2652 47354 2658 47356
rect 2412 47302 2414 47354
rect 2594 47302 2596 47354
rect 2350 47300 2356 47302
rect 2412 47300 2436 47302
rect 2492 47300 2516 47302
rect 2572 47300 2596 47302
rect 2652 47300 2658 47302
rect 2350 47291 2658 47300
rect 33070 47356 33378 47365
rect 33070 47354 33076 47356
rect 33132 47354 33156 47356
rect 33212 47354 33236 47356
rect 33292 47354 33316 47356
rect 33372 47354 33378 47356
rect 33132 47302 33134 47354
rect 33314 47302 33316 47354
rect 33070 47300 33076 47302
rect 33132 47300 33156 47302
rect 33212 47300 33236 47302
rect 33292 47300 33316 47302
rect 33372 47300 33378 47302
rect 33070 47291 33378 47300
rect 3010 46812 3318 46821
rect 3010 46810 3016 46812
rect 3072 46810 3096 46812
rect 3152 46810 3176 46812
rect 3232 46810 3256 46812
rect 3312 46810 3318 46812
rect 3072 46758 3074 46810
rect 3254 46758 3256 46810
rect 3010 46756 3016 46758
rect 3072 46756 3096 46758
rect 3152 46756 3176 46758
rect 3232 46756 3256 46758
rect 3312 46756 3318 46758
rect 3010 46747 3318 46756
rect 33730 46812 34038 46821
rect 33730 46810 33736 46812
rect 33792 46810 33816 46812
rect 33872 46810 33896 46812
rect 33952 46810 33976 46812
rect 34032 46810 34038 46812
rect 33792 46758 33794 46810
rect 33974 46758 33976 46810
rect 33730 46756 33736 46758
rect 33792 46756 33816 46758
rect 33872 46756 33896 46758
rect 33952 46756 33976 46758
rect 34032 46756 34038 46758
rect 33730 46747 34038 46756
rect 2350 46268 2658 46277
rect 2350 46266 2356 46268
rect 2412 46266 2436 46268
rect 2492 46266 2516 46268
rect 2572 46266 2596 46268
rect 2652 46266 2658 46268
rect 2412 46214 2414 46266
rect 2594 46214 2596 46266
rect 2350 46212 2356 46214
rect 2412 46212 2436 46214
rect 2492 46212 2516 46214
rect 2572 46212 2596 46214
rect 2652 46212 2658 46214
rect 2350 46203 2658 46212
rect 33070 46268 33378 46277
rect 33070 46266 33076 46268
rect 33132 46266 33156 46268
rect 33212 46266 33236 46268
rect 33292 46266 33316 46268
rect 33372 46266 33378 46268
rect 33132 46214 33134 46266
rect 33314 46214 33316 46266
rect 33070 46212 33076 46214
rect 33132 46212 33156 46214
rect 33212 46212 33236 46214
rect 33292 46212 33316 46214
rect 33372 46212 33378 46214
rect 33070 46203 33378 46212
rect 3010 45724 3318 45733
rect 3010 45722 3016 45724
rect 3072 45722 3096 45724
rect 3152 45722 3176 45724
rect 3232 45722 3256 45724
rect 3312 45722 3318 45724
rect 3072 45670 3074 45722
rect 3254 45670 3256 45722
rect 3010 45668 3016 45670
rect 3072 45668 3096 45670
rect 3152 45668 3176 45670
rect 3232 45668 3256 45670
rect 3312 45668 3318 45670
rect 3010 45659 3318 45668
rect 33730 45724 34038 45733
rect 33730 45722 33736 45724
rect 33792 45722 33816 45724
rect 33872 45722 33896 45724
rect 33952 45722 33976 45724
rect 34032 45722 34038 45724
rect 33792 45670 33794 45722
rect 33974 45670 33976 45722
rect 33730 45668 33736 45670
rect 33792 45668 33816 45670
rect 33872 45668 33896 45670
rect 33952 45668 33976 45670
rect 34032 45668 34038 45670
rect 33730 45659 34038 45668
rect 38120 45554 38148 55186
rect 38384 55208 38516 55214
rect 38436 55186 38516 55208
rect 38626 55270 38700 55298
rect 38626 55214 38654 55270
rect 40144 55214 40172 56102
rect 40236 55418 40264 56442
rect 41984 56302 42012 57394
rect 43916 56438 43944 57394
rect 43904 56432 43956 56438
rect 43904 56374 43956 56380
rect 41604 56296 41656 56302
rect 41604 56238 41656 56244
rect 41972 56296 42024 56302
rect 41972 56238 42024 56244
rect 43720 56296 43772 56302
rect 43720 56238 43772 56244
rect 41616 55418 41644 56238
rect 41972 56160 42024 56166
rect 41972 56102 42024 56108
rect 43444 56160 43496 56166
rect 43444 56102 43496 56108
rect 40224 55412 40276 55418
rect 40224 55354 40276 55360
rect 41604 55412 41656 55418
rect 41604 55354 41656 55360
rect 38626 55186 38700 55214
rect 38384 55150 38436 55156
rect 38672 55078 38700 55186
rect 40132 55208 40184 55214
rect 40132 55150 40184 55156
rect 39856 55140 39908 55146
rect 39856 55082 39908 55088
rect 38660 55072 38712 55078
rect 38660 55014 38712 55020
rect 39868 54874 39896 55082
rect 39856 54868 39908 54874
rect 39856 54810 39908 54816
rect 41984 54602 42012 56102
rect 43456 55758 43484 56102
rect 43732 55962 43760 56238
rect 43720 55956 43772 55962
rect 43720 55898 43772 55904
rect 43916 55758 43944 56374
rect 45008 56296 45060 56302
rect 45008 56238 45060 56244
rect 44364 56160 44416 56166
rect 44364 56102 44416 56108
rect 44916 56160 44968 56166
rect 44916 56102 44968 56108
rect 44376 55758 44404 56102
rect 44928 55758 44956 56102
rect 45020 55962 45048 56238
rect 45008 55956 45060 55962
rect 45008 55898 45060 55904
rect 45572 55758 45600 57394
rect 47688 56438 47716 57394
rect 49436 56506 49464 57394
rect 51080 56976 51132 56982
rect 51080 56918 51132 56924
rect 49424 56500 49476 56506
rect 49424 56442 49476 56448
rect 49792 56500 49844 56506
rect 49792 56442 49844 56448
rect 46940 56432 46992 56438
rect 46940 56374 46992 56380
rect 47676 56432 47728 56438
rect 47676 56374 47728 56380
rect 45836 56364 45888 56370
rect 45836 56306 45888 56312
rect 43444 55752 43496 55758
rect 43444 55694 43496 55700
rect 43904 55752 43956 55758
rect 43904 55694 43956 55700
rect 44364 55752 44416 55758
rect 44364 55694 44416 55700
rect 44916 55752 44968 55758
rect 44916 55694 44968 55700
rect 45560 55752 45612 55758
rect 45560 55694 45612 55700
rect 43260 55616 43312 55622
rect 43260 55558 43312 55564
rect 43272 55350 43300 55558
rect 43260 55344 43312 55350
rect 43260 55286 43312 55292
rect 42984 55208 43036 55214
rect 42984 55150 43036 55156
rect 42996 54738 43024 55150
rect 43916 54874 43944 55694
rect 44732 55684 44784 55690
rect 44732 55626 44784 55632
rect 44548 55616 44600 55622
rect 44548 55558 44600 55564
rect 44640 55616 44692 55622
rect 44640 55558 44692 55564
rect 44560 55214 44588 55558
rect 44272 55208 44324 55214
rect 44272 55150 44324 55156
rect 44548 55208 44600 55214
rect 44548 55150 44600 55156
rect 43904 54868 43956 54874
rect 43904 54810 43956 54816
rect 42984 54732 43036 54738
rect 42984 54674 43036 54680
rect 44284 54670 44312 55150
rect 44272 54664 44324 54670
rect 44272 54606 44324 54612
rect 41972 54596 42024 54602
rect 41972 54538 42024 54544
rect 44652 54262 44680 55558
rect 44744 55418 44772 55626
rect 44732 55412 44784 55418
rect 44732 55354 44784 55360
rect 45192 55208 45244 55214
rect 45192 55150 45244 55156
rect 45204 54670 45232 55150
rect 44824 54664 44876 54670
rect 44824 54606 44876 54612
rect 45192 54664 45244 54670
rect 45192 54606 45244 54612
rect 44836 54262 44864 54606
rect 44640 54256 44692 54262
rect 44640 54198 44692 54204
rect 44824 54256 44876 54262
rect 44824 54198 44876 54204
rect 45848 54126 45876 56306
rect 46756 55412 46808 55418
rect 46756 55354 46808 55360
rect 46768 55282 46796 55354
rect 46756 55276 46808 55282
rect 46756 55218 46808 55224
rect 46768 54738 46796 55218
rect 46952 55214 46980 56374
rect 49056 56296 49108 56302
rect 49056 56238 49108 56244
rect 49068 56166 49096 56238
rect 49056 56160 49108 56166
rect 49056 56102 49108 56108
rect 48596 55344 48648 55350
rect 48780 55344 48832 55350
rect 48648 55292 48780 55298
rect 49068 55321 49096 56102
rect 49608 55616 49660 55622
rect 49608 55558 49660 55564
rect 49620 55350 49648 55558
rect 49608 55344 49660 55350
rect 48596 55286 48832 55292
rect 49054 55312 49110 55321
rect 48608 55270 48820 55286
rect 49608 55286 49660 55292
rect 49054 55247 49110 55256
rect 49804 55214 49832 56442
rect 51092 56370 51120 56918
rect 51184 56438 51212 57394
rect 51540 57044 51592 57050
rect 51540 56986 51592 56992
rect 51552 56914 51580 56986
rect 52012 56914 52040 57394
rect 52276 57044 52328 57050
rect 52276 56986 52328 56992
rect 51540 56908 51592 56914
rect 51540 56850 51592 56856
rect 52000 56908 52052 56914
rect 52000 56850 52052 56856
rect 51172 56432 51224 56438
rect 51172 56374 51224 56380
rect 51080 56364 51132 56370
rect 51080 56306 51132 56312
rect 51080 56160 51132 56166
rect 51080 56102 51132 56108
rect 51092 55350 51120 56102
rect 51080 55344 51132 55350
rect 51080 55286 51132 55292
rect 51184 55214 51212 56374
rect 51552 56302 51580 56850
rect 51632 56704 51684 56710
rect 51632 56646 51684 56652
rect 51540 56296 51592 56302
rect 51540 56238 51592 56244
rect 51644 55826 51672 56646
rect 52012 56506 52040 56850
rect 52000 56500 52052 56506
rect 52000 56442 52052 56448
rect 52288 56302 52316 56986
rect 53024 56914 53052 57462
rect 55864 57452 55916 57458
rect 55864 57394 55916 57400
rect 53012 56908 53064 56914
rect 53012 56850 53064 56856
rect 52736 56840 52788 56846
rect 52736 56782 52788 56788
rect 52460 56704 52512 56710
rect 52460 56646 52512 56652
rect 52472 56370 52500 56646
rect 52748 56506 52776 56782
rect 52920 56704 52972 56710
rect 52920 56646 52972 56652
rect 52552 56500 52604 56506
rect 52552 56442 52604 56448
rect 52736 56500 52788 56506
rect 52736 56442 52788 56448
rect 52460 56364 52512 56370
rect 52460 56306 52512 56312
rect 52276 56296 52328 56302
rect 52276 56238 52328 56244
rect 51724 56228 51776 56234
rect 51724 56170 51776 56176
rect 51632 55820 51684 55826
rect 51632 55762 51684 55768
rect 51356 55752 51408 55758
rect 51356 55694 51408 55700
rect 51368 55418 51396 55694
rect 51540 55616 51592 55622
rect 51540 55558 51592 55564
rect 51356 55412 51408 55418
rect 51356 55354 51408 55360
rect 46940 55208 46992 55214
rect 46940 55150 46992 55156
rect 49792 55208 49844 55214
rect 49792 55150 49844 55156
rect 51172 55208 51224 55214
rect 51172 55150 51224 55156
rect 51368 54738 51396 55354
rect 51552 55350 51580 55558
rect 51540 55344 51592 55350
rect 51540 55286 51592 55292
rect 51736 55214 51764 56170
rect 52000 56160 52052 56166
rect 52000 56102 52052 56108
rect 51724 55208 51776 55214
rect 51724 55150 51776 55156
rect 52012 54738 52040 56102
rect 52564 55214 52592 56442
rect 52932 56438 52960 56646
rect 52920 56432 52972 56438
rect 52920 56374 52972 56380
rect 52920 55956 52972 55962
rect 52920 55898 52972 55904
rect 52644 55616 52696 55622
rect 52644 55558 52696 55564
rect 52552 55208 52604 55214
rect 52552 55150 52604 55156
rect 52656 54738 52684 55558
rect 52932 55350 52960 55898
rect 52920 55344 52972 55350
rect 52920 55286 52972 55292
rect 53024 54874 53052 56850
rect 55876 56438 55904 57394
rect 55220 56432 55272 56438
rect 55220 56374 55272 56380
rect 55864 56432 55916 56438
rect 55864 56374 55916 56380
rect 55232 55418 55260 56374
rect 56152 56370 56180 57462
rect 55312 56364 55364 56370
rect 55312 56306 55364 56312
rect 56140 56364 56192 56370
rect 56140 56306 56192 56312
rect 55324 55962 55352 56306
rect 55312 55956 55364 55962
rect 55312 55898 55364 55904
rect 55220 55412 55272 55418
rect 55220 55354 55272 55360
rect 53472 55344 53524 55350
rect 53472 55286 53524 55292
rect 53012 54868 53064 54874
rect 53012 54810 53064 54816
rect 46756 54732 46808 54738
rect 46756 54674 46808 54680
rect 51356 54732 51408 54738
rect 51356 54674 51408 54680
rect 52000 54732 52052 54738
rect 52000 54674 52052 54680
rect 52644 54732 52696 54738
rect 52644 54674 52696 54680
rect 46768 54330 46796 54674
rect 53484 54670 53512 55286
rect 53472 54664 53524 54670
rect 53472 54606 53524 54612
rect 58256 54664 58308 54670
rect 58256 54606 58308 54612
rect 46756 54324 46808 54330
rect 46756 54266 46808 54272
rect 45836 54120 45888 54126
rect 45836 54062 45888 54068
rect 38028 45526 38148 45554
rect 2350 45180 2658 45189
rect 2350 45178 2356 45180
rect 2412 45178 2436 45180
rect 2492 45178 2516 45180
rect 2572 45178 2596 45180
rect 2652 45178 2658 45180
rect 2412 45126 2414 45178
rect 2594 45126 2596 45178
rect 2350 45124 2356 45126
rect 2412 45124 2436 45126
rect 2492 45124 2516 45126
rect 2572 45124 2596 45126
rect 2652 45124 2658 45126
rect 2350 45115 2658 45124
rect 33070 45180 33378 45189
rect 33070 45178 33076 45180
rect 33132 45178 33156 45180
rect 33212 45178 33236 45180
rect 33292 45178 33316 45180
rect 33372 45178 33378 45180
rect 33132 45126 33134 45178
rect 33314 45126 33316 45178
rect 33070 45124 33076 45126
rect 33132 45124 33156 45126
rect 33212 45124 33236 45126
rect 33292 45124 33316 45126
rect 33372 45124 33378 45126
rect 33070 45115 33378 45124
rect 3010 44636 3318 44645
rect 3010 44634 3016 44636
rect 3072 44634 3096 44636
rect 3152 44634 3176 44636
rect 3232 44634 3256 44636
rect 3312 44634 3318 44636
rect 3072 44582 3074 44634
rect 3254 44582 3256 44634
rect 3010 44580 3016 44582
rect 3072 44580 3096 44582
rect 3152 44580 3176 44582
rect 3232 44580 3256 44582
rect 3312 44580 3318 44582
rect 3010 44571 3318 44580
rect 33730 44636 34038 44645
rect 33730 44634 33736 44636
rect 33792 44634 33816 44636
rect 33872 44634 33896 44636
rect 33952 44634 33976 44636
rect 34032 44634 34038 44636
rect 33792 44582 33794 44634
rect 33974 44582 33976 44634
rect 33730 44580 33736 44582
rect 33792 44580 33816 44582
rect 33872 44580 33896 44582
rect 33952 44580 33976 44582
rect 34032 44580 34038 44582
rect 33730 44571 34038 44580
rect 2350 44092 2658 44101
rect 2350 44090 2356 44092
rect 2412 44090 2436 44092
rect 2492 44090 2516 44092
rect 2572 44090 2596 44092
rect 2652 44090 2658 44092
rect 2412 44038 2414 44090
rect 2594 44038 2596 44090
rect 2350 44036 2356 44038
rect 2412 44036 2436 44038
rect 2492 44036 2516 44038
rect 2572 44036 2596 44038
rect 2652 44036 2658 44038
rect 2350 44027 2658 44036
rect 33070 44092 33378 44101
rect 33070 44090 33076 44092
rect 33132 44090 33156 44092
rect 33212 44090 33236 44092
rect 33292 44090 33316 44092
rect 33372 44090 33378 44092
rect 33132 44038 33134 44090
rect 33314 44038 33316 44090
rect 33070 44036 33076 44038
rect 33132 44036 33156 44038
rect 33212 44036 33236 44038
rect 33292 44036 33316 44038
rect 33372 44036 33378 44038
rect 33070 44027 33378 44036
rect 3010 43548 3318 43557
rect 3010 43546 3016 43548
rect 3072 43546 3096 43548
rect 3152 43546 3176 43548
rect 3232 43546 3256 43548
rect 3312 43546 3318 43548
rect 3072 43494 3074 43546
rect 3254 43494 3256 43546
rect 3010 43492 3016 43494
rect 3072 43492 3096 43494
rect 3152 43492 3176 43494
rect 3232 43492 3256 43494
rect 3312 43492 3318 43494
rect 3010 43483 3318 43492
rect 33730 43548 34038 43557
rect 33730 43546 33736 43548
rect 33792 43546 33816 43548
rect 33872 43546 33896 43548
rect 33952 43546 33976 43548
rect 34032 43546 34038 43548
rect 33792 43494 33794 43546
rect 33974 43494 33976 43546
rect 33730 43492 33736 43494
rect 33792 43492 33816 43494
rect 33872 43492 33896 43494
rect 33952 43492 33976 43494
rect 34032 43492 34038 43494
rect 33730 43483 34038 43492
rect 2350 43004 2658 43013
rect 2350 43002 2356 43004
rect 2412 43002 2436 43004
rect 2492 43002 2516 43004
rect 2572 43002 2596 43004
rect 2652 43002 2658 43004
rect 2412 42950 2414 43002
rect 2594 42950 2596 43002
rect 2350 42948 2356 42950
rect 2412 42948 2436 42950
rect 2492 42948 2516 42950
rect 2572 42948 2596 42950
rect 2652 42948 2658 42950
rect 2350 42939 2658 42948
rect 33070 43004 33378 43013
rect 33070 43002 33076 43004
rect 33132 43002 33156 43004
rect 33212 43002 33236 43004
rect 33292 43002 33316 43004
rect 33372 43002 33378 43004
rect 33132 42950 33134 43002
rect 33314 42950 33316 43002
rect 33070 42948 33076 42950
rect 33132 42948 33156 42950
rect 33212 42948 33236 42950
rect 33292 42948 33316 42950
rect 33372 42948 33378 42950
rect 33070 42939 33378 42948
rect 3010 42460 3318 42469
rect 3010 42458 3016 42460
rect 3072 42458 3096 42460
rect 3152 42458 3176 42460
rect 3232 42458 3256 42460
rect 3312 42458 3318 42460
rect 3072 42406 3074 42458
rect 3254 42406 3256 42458
rect 3010 42404 3016 42406
rect 3072 42404 3096 42406
rect 3152 42404 3176 42406
rect 3232 42404 3256 42406
rect 3312 42404 3318 42406
rect 3010 42395 3318 42404
rect 33730 42460 34038 42469
rect 33730 42458 33736 42460
rect 33792 42458 33816 42460
rect 33872 42458 33896 42460
rect 33952 42458 33976 42460
rect 34032 42458 34038 42460
rect 33792 42406 33794 42458
rect 33974 42406 33976 42458
rect 33730 42404 33736 42406
rect 33792 42404 33816 42406
rect 33872 42404 33896 42406
rect 33952 42404 33976 42406
rect 34032 42404 34038 42406
rect 33730 42395 34038 42404
rect 2350 41916 2658 41925
rect 2350 41914 2356 41916
rect 2412 41914 2436 41916
rect 2492 41914 2516 41916
rect 2572 41914 2596 41916
rect 2652 41914 2658 41916
rect 2412 41862 2414 41914
rect 2594 41862 2596 41914
rect 2350 41860 2356 41862
rect 2412 41860 2436 41862
rect 2492 41860 2516 41862
rect 2572 41860 2596 41862
rect 2652 41860 2658 41862
rect 2350 41851 2658 41860
rect 33070 41916 33378 41925
rect 33070 41914 33076 41916
rect 33132 41914 33156 41916
rect 33212 41914 33236 41916
rect 33292 41914 33316 41916
rect 33372 41914 33378 41916
rect 33132 41862 33134 41914
rect 33314 41862 33316 41914
rect 33070 41860 33076 41862
rect 33132 41860 33156 41862
rect 33212 41860 33236 41862
rect 33292 41860 33316 41862
rect 33372 41860 33378 41862
rect 33070 41851 33378 41860
rect 3010 41372 3318 41381
rect 3010 41370 3016 41372
rect 3072 41370 3096 41372
rect 3152 41370 3176 41372
rect 3232 41370 3256 41372
rect 3312 41370 3318 41372
rect 3072 41318 3074 41370
rect 3254 41318 3256 41370
rect 3010 41316 3016 41318
rect 3072 41316 3096 41318
rect 3152 41316 3176 41318
rect 3232 41316 3256 41318
rect 3312 41316 3318 41318
rect 3010 41307 3318 41316
rect 33730 41372 34038 41381
rect 33730 41370 33736 41372
rect 33792 41370 33816 41372
rect 33872 41370 33896 41372
rect 33952 41370 33976 41372
rect 34032 41370 34038 41372
rect 33792 41318 33794 41370
rect 33974 41318 33976 41370
rect 33730 41316 33736 41318
rect 33792 41316 33816 41318
rect 33872 41316 33896 41318
rect 33952 41316 33976 41318
rect 34032 41316 34038 41318
rect 33730 41307 34038 41316
rect 2350 40828 2658 40837
rect 2350 40826 2356 40828
rect 2412 40826 2436 40828
rect 2492 40826 2516 40828
rect 2572 40826 2596 40828
rect 2652 40826 2658 40828
rect 2412 40774 2414 40826
rect 2594 40774 2596 40826
rect 2350 40772 2356 40774
rect 2412 40772 2436 40774
rect 2492 40772 2516 40774
rect 2572 40772 2596 40774
rect 2652 40772 2658 40774
rect 2350 40763 2658 40772
rect 33070 40828 33378 40837
rect 33070 40826 33076 40828
rect 33132 40826 33156 40828
rect 33212 40826 33236 40828
rect 33292 40826 33316 40828
rect 33372 40826 33378 40828
rect 33132 40774 33134 40826
rect 33314 40774 33316 40826
rect 33070 40772 33076 40774
rect 33132 40772 33156 40774
rect 33212 40772 33236 40774
rect 33292 40772 33316 40774
rect 33372 40772 33378 40774
rect 33070 40763 33378 40772
rect 3010 40284 3318 40293
rect 3010 40282 3016 40284
rect 3072 40282 3096 40284
rect 3152 40282 3176 40284
rect 3232 40282 3256 40284
rect 3312 40282 3318 40284
rect 3072 40230 3074 40282
rect 3254 40230 3256 40282
rect 3010 40228 3016 40230
rect 3072 40228 3096 40230
rect 3152 40228 3176 40230
rect 3232 40228 3256 40230
rect 3312 40228 3318 40230
rect 3010 40219 3318 40228
rect 33730 40284 34038 40293
rect 33730 40282 33736 40284
rect 33792 40282 33816 40284
rect 33872 40282 33896 40284
rect 33952 40282 33976 40284
rect 34032 40282 34038 40284
rect 33792 40230 33794 40282
rect 33974 40230 33976 40282
rect 33730 40228 33736 40230
rect 33792 40228 33816 40230
rect 33872 40228 33896 40230
rect 33952 40228 33976 40230
rect 34032 40228 34038 40230
rect 33730 40219 34038 40228
rect 2350 39740 2658 39749
rect 2350 39738 2356 39740
rect 2412 39738 2436 39740
rect 2492 39738 2516 39740
rect 2572 39738 2596 39740
rect 2652 39738 2658 39740
rect 2412 39686 2414 39738
rect 2594 39686 2596 39738
rect 2350 39684 2356 39686
rect 2412 39684 2436 39686
rect 2492 39684 2516 39686
rect 2572 39684 2596 39686
rect 2652 39684 2658 39686
rect 2350 39675 2658 39684
rect 33070 39740 33378 39749
rect 33070 39738 33076 39740
rect 33132 39738 33156 39740
rect 33212 39738 33236 39740
rect 33292 39738 33316 39740
rect 33372 39738 33378 39740
rect 33132 39686 33134 39738
rect 33314 39686 33316 39738
rect 33070 39684 33076 39686
rect 33132 39684 33156 39686
rect 33212 39684 33236 39686
rect 33292 39684 33316 39686
rect 33372 39684 33378 39686
rect 33070 39675 33378 39684
rect 3010 39196 3318 39205
rect 3010 39194 3016 39196
rect 3072 39194 3096 39196
rect 3152 39194 3176 39196
rect 3232 39194 3256 39196
rect 3312 39194 3318 39196
rect 3072 39142 3074 39194
rect 3254 39142 3256 39194
rect 3010 39140 3016 39142
rect 3072 39140 3096 39142
rect 3152 39140 3176 39142
rect 3232 39140 3256 39142
rect 3312 39140 3318 39142
rect 3010 39131 3318 39140
rect 33730 39196 34038 39205
rect 33730 39194 33736 39196
rect 33792 39194 33816 39196
rect 33872 39194 33896 39196
rect 33952 39194 33976 39196
rect 34032 39194 34038 39196
rect 33792 39142 33794 39194
rect 33974 39142 33976 39194
rect 33730 39140 33736 39142
rect 33792 39140 33816 39142
rect 33872 39140 33896 39142
rect 33952 39140 33976 39142
rect 34032 39140 34038 39142
rect 33730 39131 34038 39140
rect 2350 38652 2658 38661
rect 2350 38650 2356 38652
rect 2412 38650 2436 38652
rect 2492 38650 2516 38652
rect 2572 38650 2596 38652
rect 2652 38650 2658 38652
rect 2412 38598 2414 38650
rect 2594 38598 2596 38650
rect 2350 38596 2356 38598
rect 2412 38596 2436 38598
rect 2492 38596 2516 38598
rect 2572 38596 2596 38598
rect 2652 38596 2658 38598
rect 2350 38587 2658 38596
rect 33070 38652 33378 38661
rect 33070 38650 33076 38652
rect 33132 38650 33156 38652
rect 33212 38650 33236 38652
rect 33292 38650 33316 38652
rect 33372 38650 33378 38652
rect 33132 38598 33134 38650
rect 33314 38598 33316 38650
rect 33070 38596 33076 38598
rect 33132 38596 33156 38598
rect 33212 38596 33236 38598
rect 33292 38596 33316 38598
rect 33372 38596 33378 38598
rect 33070 38587 33378 38596
rect 3010 38108 3318 38117
rect 3010 38106 3016 38108
rect 3072 38106 3096 38108
rect 3152 38106 3176 38108
rect 3232 38106 3256 38108
rect 3312 38106 3318 38108
rect 3072 38054 3074 38106
rect 3254 38054 3256 38106
rect 3010 38052 3016 38054
rect 3072 38052 3096 38054
rect 3152 38052 3176 38054
rect 3232 38052 3256 38054
rect 3312 38052 3318 38054
rect 3010 38043 3318 38052
rect 33730 38108 34038 38117
rect 33730 38106 33736 38108
rect 33792 38106 33816 38108
rect 33872 38106 33896 38108
rect 33952 38106 33976 38108
rect 34032 38106 34038 38108
rect 33792 38054 33794 38106
rect 33974 38054 33976 38106
rect 33730 38052 33736 38054
rect 33792 38052 33816 38054
rect 33872 38052 33896 38054
rect 33952 38052 33976 38054
rect 34032 38052 34038 38054
rect 33730 38043 34038 38052
rect 2350 37564 2658 37573
rect 2350 37562 2356 37564
rect 2412 37562 2436 37564
rect 2492 37562 2516 37564
rect 2572 37562 2596 37564
rect 2652 37562 2658 37564
rect 2412 37510 2414 37562
rect 2594 37510 2596 37562
rect 2350 37508 2356 37510
rect 2412 37508 2436 37510
rect 2492 37508 2516 37510
rect 2572 37508 2596 37510
rect 2652 37508 2658 37510
rect 2350 37499 2658 37508
rect 33070 37564 33378 37573
rect 33070 37562 33076 37564
rect 33132 37562 33156 37564
rect 33212 37562 33236 37564
rect 33292 37562 33316 37564
rect 33372 37562 33378 37564
rect 33132 37510 33134 37562
rect 33314 37510 33316 37562
rect 33070 37508 33076 37510
rect 33132 37508 33156 37510
rect 33212 37508 33236 37510
rect 33292 37508 33316 37510
rect 33372 37508 33378 37510
rect 33070 37499 33378 37508
rect 3010 37020 3318 37029
rect 3010 37018 3016 37020
rect 3072 37018 3096 37020
rect 3152 37018 3176 37020
rect 3232 37018 3256 37020
rect 3312 37018 3318 37020
rect 3072 36966 3074 37018
rect 3254 36966 3256 37018
rect 3010 36964 3016 36966
rect 3072 36964 3096 36966
rect 3152 36964 3176 36966
rect 3232 36964 3256 36966
rect 3312 36964 3318 36966
rect 3010 36955 3318 36964
rect 33730 37020 34038 37029
rect 33730 37018 33736 37020
rect 33792 37018 33816 37020
rect 33872 37018 33896 37020
rect 33952 37018 33976 37020
rect 34032 37018 34038 37020
rect 33792 36966 33794 37018
rect 33974 36966 33976 37018
rect 33730 36964 33736 36966
rect 33792 36964 33816 36966
rect 33872 36964 33896 36966
rect 33952 36964 33976 36966
rect 34032 36964 34038 36966
rect 33730 36955 34038 36964
rect 2350 36476 2658 36485
rect 2350 36474 2356 36476
rect 2412 36474 2436 36476
rect 2492 36474 2516 36476
rect 2572 36474 2596 36476
rect 2652 36474 2658 36476
rect 2412 36422 2414 36474
rect 2594 36422 2596 36474
rect 2350 36420 2356 36422
rect 2412 36420 2436 36422
rect 2492 36420 2516 36422
rect 2572 36420 2596 36422
rect 2652 36420 2658 36422
rect 2350 36411 2658 36420
rect 33070 36476 33378 36485
rect 33070 36474 33076 36476
rect 33132 36474 33156 36476
rect 33212 36474 33236 36476
rect 33292 36474 33316 36476
rect 33372 36474 33378 36476
rect 33132 36422 33134 36474
rect 33314 36422 33316 36474
rect 33070 36420 33076 36422
rect 33132 36420 33156 36422
rect 33212 36420 33236 36422
rect 33292 36420 33316 36422
rect 33372 36420 33378 36422
rect 33070 36411 33378 36420
rect 3010 35932 3318 35941
rect 3010 35930 3016 35932
rect 3072 35930 3096 35932
rect 3152 35930 3176 35932
rect 3232 35930 3256 35932
rect 3312 35930 3318 35932
rect 3072 35878 3074 35930
rect 3254 35878 3256 35930
rect 3010 35876 3016 35878
rect 3072 35876 3096 35878
rect 3152 35876 3176 35878
rect 3232 35876 3256 35878
rect 3312 35876 3318 35878
rect 3010 35867 3318 35876
rect 33730 35932 34038 35941
rect 33730 35930 33736 35932
rect 33792 35930 33816 35932
rect 33872 35930 33896 35932
rect 33952 35930 33976 35932
rect 34032 35930 34038 35932
rect 33792 35878 33794 35930
rect 33974 35878 33976 35930
rect 33730 35876 33736 35878
rect 33792 35876 33816 35878
rect 33872 35876 33896 35878
rect 33952 35876 33976 35878
rect 34032 35876 34038 35878
rect 33730 35867 34038 35876
rect 2350 35388 2658 35397
rect 2350 35386 2356 35388
rect 2412 35386 2436 35388
rect 2492 35386 2516 35388
rect 2572 35386 2596 35388
rect 2652 35386 2658 35388
rect 2412 35334 2414 35386
rect 2594 35334 2596 35386
rect 2350 35332 2356 35334
rect 2412 35332 2436 35334
rect 2492 35332 2516 35334
rect 2572 35332 2596 35334
rect 2652 35332 2658 35334
rect 2350 35323 2658 35332
rect 33070 35388 33378 35397
rect 33070 35386 33076 35388
rect 33132 35386 33156 35388
rect 33212 35386 33236 35388
rect 33292 35386 33316 35388
rect 33372 35386 33378 35388
rect 33132 35334 33134 35386
rect 33314 35334 33316 35386
rect 33070 35332 33076 35334
rect 33132 35332 33156 35334
rect 33212 35332 33236 35334
rect 33292 35332 33316 35334
rect 33372 35332 33378 35334
rect 33070 35323 33378 35332
rect 3010 34844 3318 34853
rect 3010 34842 3016 34844
rect 3072 34842 3096 34844
rect 3152 34842 3176 34844
rect 3232 34842 3256 34844
rect 3312 34842 3318 34844
rect 3072 34790 3074 34842
rect 3254 34790 3256 34842
rect 3010 34788 3016 34790
rect 3072 34788 3096 34790
rect 3152 34788 3176 34790
rect 3232 34788 3256 34790
rect 3312 34788 3318 34790
rect 3010 34779 3318 34788
rect 33730 34844 34038 34853
rect 33730 34842 33736 34844
rect 33792 34842 33816 34844
rect 33872 34842 33896 34844
rect 33952 34842 33976 34844
rect 34032 34842 34038 34844
rect 33792 34790 33794 34842
rect 33974 34790 33976 34842
rect 33730 34788 33736 34790
rect 33792 34788 33816 34790
rect 33872 34788 33896 34790
rect 33952 34788 33976 34790
rect 34032 34788 34038 34790
rect 33730 34779 34038 34788
rect 2350 34300 2658 34309
rect 2350 34298 2356 34300
rect 2412 34298 2436 34300
rect 2492 34298 2516 34300
rect 2572 34298 2596 34300
rect 2652 34298 2658 34300
rect 2412 34246 2414 34298
rect 2594 34246 2596 34298
rect 2350 34244 2356 34246
rect 2412 34244 2436 34246
rect 2492 34244 2516 34246
rect 2572 34244 2596 34246
rect 2652 34244 2658 34246
rect 2350 34235 2658 34244
rect 33070 34300 33378 34309
rect 33070 34298 33076 34300
rect 33132 34298 33156 34300
rect 33212 34298 33236 34300
rect 33292 34298 33316 34300
rect 33372 34298 33378 34300
rect 33132 34246 33134 34298
rect 33314 34246 33316 34298
rect 33070 34244 33076 34246
rect 33132 34244 33156 34246
rect 33212 34244 33236 34246
rect 33292 34244 33316 34246
rect 33372 34244 33378 34246
rect 33070 34235 33378 34244
rect 3010 33756 3318 33765
rect 3010 33754 3016 33756
rect 3072 33754 3096 33756
rect 3152 33754 3176 33756
rect 3232 33754 3256 33756
rect 3312 33754 3318 33756
rect 3072 33702 3074 33754
rect 3254 33702 3256 33754
rect 3010 33700 3016 33702
rect 3072 33700 3096 33702
rect 3152 33700 3176 33702
rect 3232 33700 3256 33702
rect 3312 33700 3318 33702
rect 3010 33691 3318 33700
rect 33730 33756 34038 33765
rect 33730 33754 33736 33756
rect 33792 33754 33816 33756
rect 33872 33754 33896 33756
rect 33952 33754 33976 33756
rect 34032 33754 34038 33756
rect 33792 33702 33794 33754
rect 33974 33702 33976 33754
rect 33730 33700 33736 33702
rect 33792 33700 33816 33702
rect 33872 33700 33896 33702
rect 33952 33700 33976 33702
rect 34032 33700 34038 33702
rect 33730 33691 34038 33700
rect 2350 33212 2658 33221
rect 2350 33210 2356 33212
rect 2412 33210 2436 33212
rect 2492 33210 2516 33212
rect 2572 33210 2596 33212
rect 2652 33210 2658 33212
rect 2412 33158 2414 33210
rect 2594 33158 2596 33210
rect 2350 33156 2356 33158
rect 2412 33156 2436 33158
rect 2492 33156 2516 33158
rect 2572 33156 2596 33158
rect 2652 33156 2658 33158
rect 2350 33147 2658 33156
rect 33070 33212 33378 33221
rect 33070 33210 33076 33212
rect 33132 33210 33156 33212
rect 33212 33210 33236 33212
rect 33292 33210 33316 33212
rect 33372 33210 33378 33212
rect 33132 33158 33134 33210
rect 33314 33158 33316 33210
rect 33070 33156 33076 33158
rect 33132 33156 33156 33158
rect 33212 33156 33236 33158
rect 33292 33156 33316 33158
rect 33372 33156 33378 33158
rect 33070 33147 33378 33156
rect 3010 32668 3318 32677
rect 3010 32666 3016 32668
rect 3072 32666 3096 32668
rect 3152 32666 3176 32668
rect 3232 32666 3256 32668
rect 3312 32666 3318 32668
rect 3072 32614 3074 32666
rect 3254 32614 3256 32666
rect 3010 32612 3016 32614
rect 3072 32612 3096 32614
rect 3152 32612 3176 32614
rect 3232 32612 3256 32614
rect 3312 32612 3318 32614
rect 3010 32603 3318 32612
rect 33730 32668 34038 32677
rect 33730 32666 33736 32668
rect 33792 32666 33816 32668
rect 33872 32666 33896 32668
rect 33952 32666 33976 32668
rect 34032 32666 34038 32668
rect 33792 32614 33794 32666
rect 33974 32614 33976 32666
rect 33730 32612 33736 32614
rect 33792 32612 33816 32614
rect 33872 32612 33896 32614
rect 33952 32612 33976 32614
rect 34032 32612 34038 32614
rect 33730 32603 34038 32612
rect 2350 32124 2658 32133
rect 2350 32122 2356 32124
rect 2412 32122 2436 32124
rect 2492 32122 2516 32124
rect 2572 32122 2596 32124
rect 2652 32122 2658 32124
rect 2412 32070 2414 32122
rect 2594 32070 2596 32122
rect 2350 32068 2356 32070
rect 2412 32068 2436 32070
rect 2492 32068 2516 32070
rect 2572 32068 2596 32070
rect 2652 32068 2658 32070
rect 2350 32059 2658 32068
rect 33070 32124 33378 32133
rect 33070 32122 33076 32124
rect 33132 32122 33156 32124
rect 33212 32122 33236 32124
rect 33292 32122 33316 32124
rect 33372 32122 33378 32124
rect 33132 32070 33134 32122
rect 33314 32070 33316 32122
rect 33070 32068 33076 32070
rect 33132 32068 33156 32070
rect 33212 32068 33236 32070
rect 33292 32068 33316 32070
rect 33372 32068 33378 32070
rect 33070 32059 33378 32068
rect 3010 31580 3318 31589
rect 3010 31578 3016 31580
rect 3072 31578 3096 31580
rect 3152 31578 3176 31580
rect 3232 31578 3256 31580
rect 3312 31578 3318 31580
rect 3072 31526 3074 31578
rect 3254 31526 3256 31578
rect 3010 31524 3016 31526
rect 3072 31524 3096 31526
rect 3152 31524 3176 31526
rect 3232 31524 3256 31526
rect 3312 31524 3318 31526
rect 3010 31515 3318 31524
rect 33730 31580 34038 31589
rect 33730 31578 33736 31580
rect 33792 31578 33816 31580
rect 33872 31578 33896 31580
rect 33952 31578 33976 31580
rect 34032 31578 34038 31580
rect 33792 31526 33794 31578
rect 33974 31526 33976 31578
rect 33730 31524 33736 31526
rect 33792 31524 33816 31526
rect 33872 31524 33896 31526
rect 33952 31524 33976 31526
rect 34032 31524 34038 31526
rect 33730 31515 34038 31524
rect 2350 31036 2658 31045
rect 2350 31034 2356 31036
rect 2412 31034 2436 31036
rect 2492 31034 2516 31036
rect 2572 31034 2596 31036
rect 2652 31034 2658 31036
rect 2412 30982 2414 31034
rect 2594 30982 2596 31034
rect 2350 30980 2356 30982
rect 2412 30980 2436 30982
rect 2492 30980 2516 30982
rect 2572 30980 2596 30982
rect 2652 30980 2658 30982
rect 2350 30971 2658 30980
rect 33070 31036 33378 31045
rect 33070 31034 33076 31036
rect 33132 31034 33156 31036
rect 33212 31034 33236 31036
rect 33292 31034 33316 31036
rect 33372 31034 33378 31036
rect 33132 30982 33134 31034
rect 33314 30982 33316 31034
rect 33070 30980 33076 30982
rect 33132 30980 33156 30982
rect 33212 30980 33236 30982
rect 33292 30980 33316 30982
rect 33372 30980 33378 30982
rect 33070 30971 33378 30980
rect 3010 30492 3318 30501
rect 3010 30490 3016 30492
rect 3072 30490 3096 30492
rect 3152 30490 3176 30492
rect 3232 30490 3256 30492
rect 3312 30490 3318 30492
rect 3072 30438 3074 30490
rect 3254 30438 3256 30490
rect 3010 30436 3016 30438
rect 3072 30436 3096 30438
rect 3152 30436 3176 30438
rect 3232 30436 3256 30438
rect 3312 30436 3318 30438
rect 3010 30427 3318 30436
rect 33730 30492 34038 30501
rect 33730 30490 33736 30492
rect 33792 30490 33816 30492
rect 33872 30490 33896 30492
rect 33952 30490 33976 30492
rect 34032 30490 34038 30492
rect 33792 30438 33794 30490
rect 33974 30438 33976 30490
rect 33730 30436 33736 30438
rect 33792 30436 33816 30438
rect 33872 30436 33896 30438
rect 33952 30436 33976 30438
rect 34032 30436 34038 30438
rect 33730 30427 34038 30436
rect 2350 29948 2658 29957
rect 2350 29946 2356 29948
rect 2412 29946 2436 29948
rect 2492 29946 2516 29948
rect 2572 29946 2596 29948
rect 2652 29946 2658 29948
rect 2412 29894 2414 29946
rect 2594 29894 2596 29946
rect 2350 29892 2356 29894
rect 2412 29892 2436 29894
rect 2492 29892 2516 29894
rect 2572 29892 2596 29894
rect 2652 29892 2658 29894
rect 2350 29883 2658 29892
rect 33070 29948 33378 29957
rect 33070 29946 33076 29948
rect 33132 29946 33156 29948
rect 33212 29946 33236 29948
rect 33292 29946 33316 29948
rect 33372 29946 33378 29948
rect 33132 29894 33134 29946
rect 33314 29894 33316 29946
rect 33070 29892 33076 29894
rect 33132 29892 33156 29894
rect 33212 29892 33236 29894
rect 33292 29892 33316 29894
rect 33372 29892 33378 29894
rect 33070 29883 33378 29892
rect 3010 29404 3318 29413
rect 3010 29402 3016 29404
rect 3072 29402 3096 29404
rect 3152 29402 3176 29404
rect 3232 29402 3256 29404
rect 3312 29402 3318 29404
rect 3072 29350 3074 29402
rect 3254 29350 3256 29402
rect 3010 29348 3016 29350
rect 3072 29348 3096 29350
rect 3152 29348 3176 29350
rect 3232 29348 3256 29350
rect 3312 29348 3318 29350
rect 3010 29339 3318 29348
rect 33730 29404 34038 29413
rect 33730 29402 33736 29404
rect 33792 29402 33816 29404
rect 33872 29402 33896 29404
rect 33952 29402 33976 29404
rect 34032 29402 34038 29404
rect 33792 29350 33794 29402
rect 33974 29350 33976 29402
rect 33730 29348 33736 29350
rect 33792 29348 33816 29350
rect 33872 29348 33896 29350
rect 33952 29348 33976 29350
rect 34032 29348 34038 29350
rect 33730 29339 34038 29348
rect 2350 28860 2658 28869
rect 2350 28858 2356 28860
rect 2412 28858 2436 28860
rect 2492 28858 2516 28860
rect 2572 28858 2596 28860
rect 2652 28858 2658 28860
rect 2412 28806 2414 28858
rect 2594 28806 2596 28858
rect 2350 28804 2356 28806
rect 2412 28804 2436 28806
rect 2492 28804 2516 28806
rect 2572 28804 2596 28806
rect 2652 28804 2658 28806
rect 2350 28795 2658 28804
rect 33070 28860 33378 28869
rect 33070 28858 33076 28860
rect 33132 28858 33156 28860
rect 33212 28858 33236 28860
rect 33292 28858 33316 28860
rect 33372 28858 33378 28860
rect 33132 28806 33134 28858
rect 33314 28806 33316 28858
rect 33070 28804 33076 28806
rect 33132 28804 33156 28806
rect 33212 28804 33236 28806
rect 33292 28804 33316 28806
rect 33372 28804 33378 28806
rect 33070 28795 33378 28804
rect 3010 28316 3318 28325
rect 3010 28314 3016 28316
rect 3072 28314 3096 28316
rect 3152 28314 3176 28316
rect 3232 28314 3256 28316
rect 3312 28314 3318 28316
rect 3072 28262 3074 28314
rect 3254 28262 3256 28314
rect 3010 28260 3016 28262
rect 3072 28260 3096 28262
rect 3152 28260 3176 28262
rect 3232 28260 3256 28262
rect 3312 28260 3318 28262
rect 3010 28251 3318 28260
rect 33730 28316 34038 28325
rect 33730 28314 33736 28316
rect 33792 28314 33816 28316
rect 33872 28314 33896 28316
rect 33952 28314 33976 28316
rect 34032 28314 34038 28316
rect 33792 28262 33794 28314
rect 33974 28262 33976 28314
rect 33730 28260 33736 28262
rect 33792 28260 33816 28262
rect 33872 28260 33896 28262
rect 33952 28260 33976 28262
rect 34032 28260 34038 28262
rect 33730 28251 34038 28260
rect 2350 27772 2658 27781
rect 2350 27770 2356 27772
rect 2412 27770 2436 27772
rect 2492 27770 2516 27772
rect 2572 27770 2596 27772
rect 2652 27770 2658 27772
rect 2412 27718 2414 27770
rect 2594 27718 2596 27770
rect 2350 27716 2356 27718
rect 2412 27716 2436 27718
rect 2492 27716 2516 27718
rect 2572 27716 2596 27718
rect 2652 27716 2658 27718
rect 2350 27707 2658 27716
rect 33070 27772 33378 27781
rect 33070 27770 33076 27772
rect 33132 27770 33156 27772
rect 33212 27770 33236 27772
rect 33292 27770 33316 27772
rect 33372 27770 33378 27772
rect 33132 27718 33134 27770
rect 33314 27718 33316 27770
rect 33070 27716 33076 27718
rect 33132 27716 33156 27718
rect 33212 27716 33236 27718
rect 33292 27716 33316 27718
rect 33372 27716 33378 27718
rect 33070 27707 33378 27716
rect 3010 27228 3318 27237
rect 3010 27226 3016 27228
rect 3072 27226 3096 27228
rect 3152 27226 3176 27228
rect 3232 27226 3256 27228
rect 3312 27226 3318 27228
rect 3072 27174 3074 27226
rect 3254 27174 3256 27226
rect 3010 27172 3016 27174
rect 3072 27172 3096 27174
rect 3152 27172 3176 27174
rect 3232 27172 3256 27174
rect 3312 27172 3318 27174
rect 3010 27163 3318 27172
rect 33730 27228 34038 27237
rect 33730 27226 33736 27228
rect 33792 27226 33816 27228
rect 33872 27226 33896 27228
rect 33952 27226 33976 27228
rect 34032 27226 34038 27228
rect 33792 27174 33794 27226
rect 33974 27174 33976 27226
rect 33730 27172 33736 27174
rect 33792 27172 33816 27174
rect 33872 27172 33896 27174
rect 33952 27172 33976 27174
rect 34032 27172 34038 27174
rect 33730 27163 34038 27172
rect 2350 26684 2658 26693
rect 2350 26682 2356 26684
rect 2412 26682 2436 26684
rect 2492 26682 2516 26684
rect 2572 26682 2596 26684
rect 2652 26682 2658 26684
rect 2412 26630 2414 26682
rect 2594 26630 2596 26682
rect 2350 26628 2356 26630
rect 2412 26628 2436 26630
rect 2492 26628 2516 26630
rect 2572 26628 2596 26630
rect 2652 26628 2658 26630
rect 2350 26619 2658 26628
rect 33070 26684 33378 26693
rect 33070 26682 33076 26684
rect 33132 26682 33156 26684
rect 33212 26682 33236 26684
rect 33292 26682 33316 26684
rect 33372 26682 33378 26684
rect 33132 26630 33134 26682
rect 33314 26630 33316 26682
rect 33070 26628 33076 26630
rect 33132 26628 33156 26630
rect 33212 26628 33236 26630
rect 33292 26628 33316 26630
rect 33372 26628 33378 26630
rect 33070 26619 33378 26628
rect 3010 26140 3318 26149
rect 3010 26138 3016 26140
rect 3072 26138 3096 26140
rect 3152 26138 3176 26140
rect 3232 26138 3256 26140
rect 3312 26138 3318 26140
rect 3072 26086 3074 26138
rect 3254 26086 3256 26138
rect 3010 26084 3016 26086
rect 3072 26084 3096 26086
rect 3152 26084 3176 26086
rect 3232 26084 3256 26086
rect 3312 26084 3318 26086
rect 3010 26075 3318 26084
rect 33730 26140 34038 26149
rect 33730 26138 33736 26140
rect 33792 26138 33816 26140
rect 33872 26138 33896 26140
rect 33952 26138 33976 26140
rect 34032 26138 34038 26140
rect 33792 26086 33794 26138
rect 33974 26086 33976 26138
rect 33730 26084 33736 26086
rect 33792 26084 33816 26086
rect 33872 26084 33896 26086
rect 33952 26084 33976 26086
rect 34032 26084 34038 26086
rect 33730 26075 34038 26084
rect 2350 25596 2658 25605
rect 2350 25594 2356 25596
rect 2412 25594 2436 25596
rect 2492 25594 2516 25596
rect 2572 25594 2596 25596
rect 2652 25594 2658 25596
rect 2412 25542 2414 25594
rect 2594 25542 2596 25594
rect 2350 25540 2356 25542
rect 2412 25540 2436 25542
rect 2492 25540 2516 25542
rect 2572 25540 2596 25542
rect 2652 25540 2658 25542
rect 2350 25531 2658 25540
rect 33070 25596 33378 25605
rect 33070 25594 33076 25596
rect 33132 25594 33156 25596
rect 33212 25594 33236 25596
rect 33292 25594 33316 25596
rect 33372 25594 33378 25596
rect 33132 25542 33134 25594
rect 33314 25542 33316 25594
rect 33070 25540 33076 25542
rect 33132 25540 33156 25542
rect 33212 25540 33236 25542
rect 33292 25540 33316 25542
rect 33372 25540 33378 25542
rect 33070 25531 33378 25540
rect 3010 25052 3318 25061
rect 3010 25050 3016 25052
rect 3072 25050 3096 25052
rect 3152 25050 3176 25052
rect 3232 25050 3256 25052
rect 3312 25050 3318 25052
rect 3072 24998 3074 25050
rect 3254 24998 3256 25050
rect 3010 24996 3016 24998
rect 3072 24996 3096 24998
rect 3152 24996 3176 24998
rect 3232 24996 3256 24998
rect 3312 24996 3318 24998
rect 3010 24987 3318 24996
rect 33730 25052 34038 25061
rect 33730 25050 33736 25052
rect 33792 25050 33816 25052
rect 33872 25050 33896 25052
rect 33952 25050 33976 25052
rect 34032 25050 34038 25052
rect 33792 24998 33794 25050
rect 33974 24998 33976 25050
rect 33730 24996 33736 24998
rect 33792 24996 33816 24998
rect 33872 24996 33896 24998
rect 33952 24996 33976 24998
rect 34032 24996 34038 24998
rect 33730 24987 34038 24996
rect 2350 24508 2658 24517
rect 2350 24506 2356 24508
rect 2412 24506 2436 24508
rect 2492 24506 2516 24508
rect 2572 24506 2596 24508
rect 2652 24506 2658 24508
rect 2412 24454 2414 24506
rect 2594 24454 2596 24506
rect 2350 24452 2356 24454
rect 2412 24452 2436 24454
rect 2492 24452 2516 24454
rect 2572 24452 2596 24454
rect 2652 24452 2658 24454
rect 2350 24443 2658 24452
rect 33070 24508 33378 24517
rect 33070 24506 33076 24508
rect 33132 24506 33156 24508
rect 33212 24506 33236 24508
rect 33292 24506 33316 24508
rect 33372 24506 33378 24508
rect 33132 24454 33134 24506
rect 33314 24454 33316 24506
rect 33070 24452 33076 24454
rect 33132 24452 33156 24454
rect 33212 24452 33236 24454
rect 33292 24452 33316 24454
rect 33372 24452 33378 24454
rect 33070 24443 33378 24452
rect 3010 23964 3318 23973
rect 3010 23962 3016 23964
rect 3072 23962 3096 23964
rect 3152 23962 3176 23964
rect 3232 23962 3256 23964
rect 3312 23962 3318 23964
rect 3072 23910 3074 23962
rect 3254 23910 3256 23962
rect 3010 23908 3016 23910
rect 3072 23908 3096 23910
rect 3152 23908 3176 23910
rect 3232 23908 3256 23910
rect 3312 23908 3318 23910
rect 3010 23899 3318 23908
rect 33730 23964 34038 23973
rect 33730 23962 33736 23964
rect 33792 23962 33816 23964
rect 33872 23962 33896 23964
rect 33952 23962 33976 23964
rect 34032 23962 34038 23964
rect 33792 23910 33794 23962
rect 33974 23910 33976 23962
rect 33730 23908 33736 23910
rect 33792 23908 33816 23910
rect 33872 23908 33896 23910
rect 33952 23908 33976 23910
rect 34032 23908 34038 23910
rect 33730 23899 34038 23908
rect 2350 23420 2658 23429
rect 2350 23418 2356 23420
rect 2412 23418 2436 23420
rect 2492 23418 2516 23420
rect 2572 23418 2596 23420
rect 2652 23418 2658 23420
rect 2412 23366 2414 23418
rect 2594 23366 2596 23418
rect 2350 23364 2356 23366
rect 2412 23364 2436 23366
rect 2492 23364 2516 23366
rect 2572 23364 2596 23366
rect 2652 23364 2658 23366
rect 2350 23355 2658 23364
rect 33070 23420 33378 23429
rect 33070 23418 33076 23420
rect 33132 23418 33156 23420
rect 33212 23418 33236 23420
rect 33292 23418 33316 23420
rect 33372 23418 33378 23420
rect 33132 23366 33134 23418
rect 33314 23366 33316 23418
rect 33070 23364 33076 23366
rect 33132 23364 33156 23366
rect 33212 23364 33236 23366
rect 33292 23364 33316 23366
rect 33372 23364 33378 23366
rect 33070 23355 33378 23364
rect 3010 22876 3318 22885
rect 3010 22874 3016 22876
rect 3072 22874 3096 22876
rect 3152 22874 3176 22876
rect 3232 22874 3256 22876
rect 3312 22874 3318 22876
rect 3072 22822 3074 22874
rect 3254 22822 3256 22874
rect 3010 22820 3016 22822
rect 3072 22820 3096 22822
rect 3152 22820 3176 22822
rect 3232 22820 3256 22822
rect 3312 22820 3318 22822
rect 3010 22811 3318 22820
rect 33730 22876 34038 22885
rect 33730 22874 33736 22876
rect 33792 22874 33816 22876
rect 33872 22874 33896 22876
rect 33952 22874 33976 22876
rect 34032 22874 34038 22876
rect 33792 22822 33794 22874
rect 33974 22822 33976 22874
rect 33730 22820 33736 22822
rect 33792 22820 33816 22822
rect 33872 22820 33896 22822
rect 33952 22820 33976 22822
rect 34032 22820 34038 22822
rect 33730 22811 34038 22820
rect 2350 22332 2658 22341
rect 2350 22330 2356 22332
rect 2412 22330 2436 22332
rect 2492 22330 2516 22332
rect 2572 22330 2596 22332
rect 2652 22330 2658 22332
rect 2412 22278 2414 22330
rect 2594 22278 2596 22330
rect 2350 22276 2356 22278
rect 2412 22276 2436 22278
rect 2492 22276 2516 22278
rect 2572 22276 2596 22278
rect 2652 22276 2658 22278
rect 2350 22267 2658 22276
rect 33070 22332 33378 22341
rect 33070 22330 33076 22332
rect 33132 22330 33156 22332
rect 33212 22330 33236 22332
rect 33292 22330 33316 22332
rect 33372 22330 33378 22332
rect 33132 22278 33134 22330
rect 33314 22278 33316 22330
rect 33070 22276 33076 22278
rect 33132 22276 33156 22278
rect 33212 22276 33236 22278
rect 33292 22276 33316 22278
rect 33372 22276 33378 22278
rect 33070 22267 33378 22276
rect 3010 21788 3318 21797
rect 3010 21786 3016 21788
rect 3072 21786 3096 21788
rect 3152 21786 3176 21788
rect 3232 21786 3256 21788
rect 3312 21786 3318 21788
rect 3072 21734 3074 21786
rect 3254 21734 3256 21786
rect 3010 21732 3016 21734
rect 3072 21732 3096 21734
rect 3152 21732 3176 21734
rect 3232 21732 3256 21734
rect 3312 21732 3318 21734
rect 3010 21723 3318 21732
rect 33730 21788 34038 21797
rect 33730 21786 33736 21788
rect 33792 21786 33816 21788
rect 33872 21786 33896 21788
rect 33952 21786 33976 21788
rect 34032 21786 34038 21788
rect 33792 21734 33794 21786
rect 33974 21734 33976 21786
rect 33730 21732 33736 21734
rect 33792 21732 33816 21734
rect 33872 21732 33896 21734
rect 33952 21732 33976 21734
rect 34032 21732 34038 21734
rect 33730 21723 34038 21732
rect 2350 21244 2658 21253
rect 2350 21242 2356 21244
rect 2412 21242 2436 21244
rect 2492 21242 2516 21244
rect 2572 21242 2596 21244
rect 2652 21242 2658 21244
rect 2412 21190 2414 21242
rect 2594 21190 2596 21242
rect 2350 21188 2356 21190
rect 2412 21188 2436 21190
rect 2492 21188 2516 21190
rect 2572 21188 2596 21190
rect 2652 21188 2658 21190
rect 2350 21179 2658 21188
rect 33070 21244 33378 21253
rect 33070 21242 33076 21244
rect 33132 21242 33156 21244
rect 33212 21242 33236 21244
rect 33292 21242 33316 21244
rect 33372 21242 33378 21244
rect 33132 21190 33134 21242
rect 33314 21190 33316 21242
rect 33070 21188 33076 21190
rect 33132 21188 33156 21190
rect 33212 21188 33236 21190
rect 33292 21188 33316 21190
rect 33372 21188 33378 21190
rect 33070 21179 33378 21188
rect 3010 20700 3318 20709
rect 3010 20698 3016 20700
rect 3072 20698 3096 20700
rect 3152 20698 3176 20700
rect 3232 20698 3256 20700
rect 3312 20698 3318 20700
rect 3072 20646 3074 20698
rect 3254 20646 3256 20698
rect 3010 20644 3016 20646
rect 3072 20644 3096 20646
rect 3152 20644 3176 20646
rect 3232 20644 3256 20646
rect 3312 20644 3318 20646
rect 3010 20635 3318 20644
rect 33730 20700 34038 20709
rect 33730 20698 33736 20700
rect 33792 20698 33816 20700
rect 33872 20698 33896 20700
rect 33952 20698 33976 20700
rect 34032 20698 34038 20700
rect 33792 20646 33794 20698
rect 33974 20646 33976 20698
rect 33730 20644 33736 20646
rect 33792 20644 33816 20646
rect 33872 20644 33896 20646
rect 33952 20644 33976 20646
rect 34032 20644 34038 20646
rect 33730 20635 34038 20644
rect 2350 20156 2658 20165
rect 2350 20154 2356 20156
rect 2412 20154 2436 20156
rect 2492 20154 2516 20156
rect 2572 20154 2596 20156
rect 2652 20154 2658 20156
rect 2412 20102 2414 20154
rect 2594 20102 2596 20154
rect 2350 20100 2356 20102
rect 2412 20100 2436 20102
rect 2492 20100 2516 20102
rect 2572 20100 2596 20102
rect 2652 20100 2658 20102
rect 2350 20091 2658 20100
rect 33070 20156 33378 20165
rect 33070 20154 33076 20156
rect 33132 20154 33156 20156
rect 33212 20154 33236 20156
rect 33292 20154 33316 20156
rect 33372 20154 33378 20156
rect 33132 20102 33134 20154
rect 33314 20102 33316 20154
rect 33070 20100 33076 20102
rect 33132 20100 33156 20102
rect 33212 20100 33236 20102
rect 33292 20100 33316 20102
rect 33372 20100 33378 20102
rect 33070 20091 33378 20100
rect 3010 19612 3318 19621
rect 3010 19610 3016 19612
rect 3072 19610 3096 19612
rect 3152 19610 3176 19612
rect 3232 19610 3256 19612
rect 3312 19610 3318 19612
rect 3072 19558 3074 19610
rect 3254 19558 3256 19610
rect 3010 19556 3016 19558
rect 3072 19556 3096 19558
rect 3152 19556 3176 19558
rect 3232 19556 3256 19558
rect 3312 19556 3318 19558
rect 3010 19547 3318 19556
rect 33730 19612 34038 19621
rect 33730 19610 33736 19612
rect 33792 19610 33816 19612
rect 33872 19610 33896 19612
rect 33952 19610 33976 19612
rect 34032 19610 34038 19612
rect 33792 19558 33794 19610
rect 33974 19558 33976 19610
rect 33730 19556 33736 19558
rect 33792 19556 33816 19558
rect 33872 19556 33896 19558
rect 33952 19556 33976 19558
rect 34032 19556 34038 19558
rect 33730 19547 34038 19556
rect 2350 19068 2658 19077
rect 2350 19066 2356 19068
rect 2412 19066 2436 19068
rect 2492 19066 2516 19068
rect 2572 19066 2596 19068
rect 2652 19066 2658 19068
rect 2412 19014 2414 19066
rect 2594 19014 2596 19066
rect 2350 19012 2356 19014
rect 2412 19012 2436 19014
rect 2492 19012 2516 19014
rect 2572 19012 2596 19014
rect 2652 19012 2658 19014
rect 2350 19003 2658 19012
rect 33070 19068 33378 19077
rect 33070 19066 33076 19068
rect 33132 19066 33156 19068
rect 33212 19066 33236 19068
rect 33292 19066 33316 19068
rect 33372 19066 33378 19068
rect 33132 19014 33134 19066
rect 33314 19014 33316 19066
rect 33070 19012 33076 19014
rect 33132 19012 33156 19014
rect 33212 19012 33236 19014
rect 33292 19012 33316 19014
rect 33372 19012 33378 19014
rect 33070 19003 33378 19012
rect 3010 18524 3318 18533
rect 3010 18522 3016 18524
rect 3072 18522 3096 18524
rect 3152 18522 3176 18524
rect 3232 18522 3256 18524
rect 3312 18522 3318 18524
rect 3072 18470 3074 18522
rect 3254 18470 3256 18522
rect 3010 18468 3016 18470
rect 3072 18468 3096 18470
rect 3152 18468 3176 18470
rect 3232 18468 3256 18470
rect 3312 18468 3318 18470
rect 3010 18459 3318 18468
rect 33730 18524 34038 18533
rect 33730 18522 33736 18524
rect 33792 18522 33816 18524
rect 33872 18522 33896 18524
rect 33952 18522 33976 18524
rect 34032 18522 34038 18524
rect 33792 18470 33794 18522
rect 33974 18470 33976 18522
rect 33730 18468 33736 18470
rect 33792 18468 33816 18470
rect 33872 18468 33896 18470
rect 33952 18468 33976 18470
rect 34032 18468 34038 18470
rect 33730 18459 34038 18468
rect 2350 17980 2658 17989
rect 2350 17978 2356 17980
rect 2412 17978 2436 17980
rect 2492 17978 2516 17980
rect 2572 17978 2596 17980
rect 2652 17978 2658 17980
rect 2412 17926 2414 17978
rect 2594 17926 2596 17978
rect 2350 17924 2356 17926
rect 2412 17924 2436 17926
rect 2492 17924 2516 17926
rect 2572 17924 2596 17926
rect 2652 17924 2658 17926
rect 2350 17915 2658 17924
rect 33070 17980 33378 17989
rect 33070 17978 33076 17980
rect 33132 17978 33156 17980
rect 33212 17978 33236 17980
rect 33292 17978 33316 17980
rect 33372 17978 33378 17980
rect 33132 17926 33134 17978
rect 33314 17926 33316 17978
rect 33070 17924 33076 17926
rect 33132 17924 33156 17926
rect 33212 17924 33236 17926
rect 33292 17924 33316 17926
rect 33372 17924 33378 17926
rect 33070 17915 33378 17924
rect 3010 17436 3318 17445
rect 3010 17434 3016 17436
rect 3072 17434 3096 17436
rect 3152 17434 3176 17436
rect 3232 17434 3256 17436
rect 3312 17434 3318 17436
rect 3072 17382 3074 17434
rect 3254 17382 3256 17434
rect 3010 17380 3016 17382
rect 3072 17380 3096 17382
rect 3152 17380 3176 17382
rect 3232 17380 3256 17382
rect 3312 17380 3318 17382
rect 3010 17371 3318 17380
rect 33730 17436 34038 17445
rect 33730 17434 33736 17436
rect 33792 17434 33816 17436
rect 33872 17434 33896 17436
rect 33952 17434 33976 17436
rect 34032 17434 34038 17436
rect 33792 17382 33794 17434
rect 33974 17382 33976 17434
rect 33730 17380 33736 17382
rect 33792 17380 33816 17382
rect 33872 17380 33896 17382
rect 33952 17380 33976 17382
rect 34032 17380 34038 17382
rect 33730 17371 34038 17380
rect 2350 16892 2658 16901
rect 2350 16890 2356 16892
rect 2412 16890 2436 16892
rect 2492 16890 2516 16892
rect 2572 16890 2596 16892
rect 2652 16890 2658 16892
rect 2412 16838 2414 16890
rect 2594 16838 2596 16890
rect 2350 16836 2356 16838
rect 2412 16836 2436 16838
rect 2492 16836 2516 16838
rect 2572 16836 2596 16838
rect 2652 16836 2658 16838
rect 2350 16827 2658 16836
rect 33070 16892 33378 16901
rect 33070 16890 33076 16892
rect 33132 16890 33156 16892
rect 33212 16890 33236 16892
rect 33292 16890 33316 16892
rect 33372 16890 33378 16892
rect 33132 16838 33134 16890
rect 33314 16838 33316 16890
rect 33070 16836 33076 16838
rect 33132 16836 33156 16838
rect 33212 16836 33236 16838
rect 33292 16836 33316 16838
rect 33372 16836 33378 16838
rect 33070 16827 33378 16836
rect 3010 16348 3318 16357
rect 3010 16346 3016 16348
rect 3072 16346 3096 16348
rect 3152 16346 3176 16348
rect 3232 16346 3256 16348
rect 3312 16346 3318 16348
rect 3072 16294 3074 16346
rect 3254 16294 3256 16346
rect 3010 16292 3016 16294
rect 3072 16292 3096 16294
rect 3152 16292 3176 16294
rect 3232 16292 3256 16294
rect 3312 16292 3318 16294
rect 3010 16283 3318 16292
rect 33730 16348 34038 16357
rect 33730 16346 33736 16348
rect 33792 16346 33816 16348
rect 33872 16346 33896 16348
rect 33952 16346 33976 16348
rect 34032 16346 34038 16348
rect 33792 16294 33794 16346
rect 33974 16294 33976 16346
rect 33730 16292 33736 16294
rect 33792 16292 33816 16294
rect 33872 16292 33896 16294
rect 33952 16292 33976 16294
rect 34032 16292 34038 16294
rect 33730 16283 34038 16292
rect 2350 15804 2658 15813
rect 2350 15802 2356 15804
rect 2412 15802 2436 15804
rect 2492 15802 2516 15804
rect 2572 15802 2596 15804
rect 2652 15802 2658 15804
rect 2412 15750 2414 15802
rect 2594 15750 2596 15802
rect 2350 15748 2356 15750
rect 2412 15748 2436 15750
rect 2492 15748 2516 15750
rect 2572 15748 2596 15750
rect 2652 15748 2658 15750
rect 2350 15739 2658 15748
rect 33070 15804 33378 15813
rect 33070 15802 33076 15804
rect 33132 15802 33156 15804
rect 33212 15802 33236 15804
rect 33292 15802 33316 15804
rect 33372 15802 33378 15804
rect 33132 15750 33134 15802
rect 33314 15750 33316 15802
rect 33070 15748 33076 15750
rect 33132 15748 33156 15750
rect 33212 15748 33236 15750
rect 33292 15748 33316 15750
rect 33372 15748 33378 15750
rect 33070 15739 33378 15748
rect 3010 15260 3318 15269
rect 3010 15258 3016 15260
rect 3072 15258 3096 15260
rect 3152 15258 3176 15260
rect 3232 15258 3256 15260
rect 3312 15258 3318 15260
rect 3072 15206 3074 15258
rect 3254 15206 3256 15258
rect 3010 15204 3016 15206
rect 3072 15204 3096 15206
rect 3152 15204 3176 15206
rect 3232 15204 3256 15206
rect 3312 15204 3318 15206
rect 3010 15195 3318 15204
rect 33730 15260 34038 15269
rect 33730 15258 33736 15260
rect 33792 15258 33816 15260
rect 33872 15258 33896 15260
rect 33952 15258 33976 15260
rect 34032 15258 34038 15260
rect 33792 15206 33794 15258
rect 33974 15206 33976 15258
rect 33730 15204 33736 15206
rect 33792 15204 33816 15206
rect 33872 15204 33896 15206
rect 33952 15204 33976 15206
rect 34032 15204 34038 15206
rect 33730 15195 34038 15204
rect 38028 15162 38056 45526
rect 58268 44946 58296 54606
rect 58530 44976 58586 44985
rect 58256 44940 58308 44946
rect 58530 44911 58586 44920
rect 58256 44882 58308 44888
rect 58544 44878 58572 44911
rect 58532 44872 58584 44878
rect 58532 44814 58584 44820
rect 38016 15156 38068 15162
rect 38016 15098 38068 15104
rect 56508 15156 56560 15162
rect 56508 15098 56560 15104
rect 56520 15065 56548 15098
rect 56506 15056 56562 15065
rect 56506 14991 56562 15000
rect 2350 14716 2658 14725
rect 2350 14714 2356 14716
rect 2412 14714 2436 14716
rect 2492 14714 2516 14716
rect 2572 14714 2596 14716
rect 2652 14714 2658 14716
rect 2412 14662 2414 14714
rect 2594 14662 2596 14714
rect 2350 14660 2356 14662
rect 2412 14660 2436 14662
rect 2492 14660 2516 14662
rect 2572 14660 2596 14662
rect 2652 14660 2658 14662
rect 2350 14651 2658 14660
rect 33070 14716 33378 14725
rect 33070 14714 33076 14716
rect 33132 14714 33156 14716
rect 33212 14714 33236 14716
rect 33292 14714 33316 14716
rect 33372 14714 33378 14716
rect 33132 14662 33134 14714
rect 33314 14662 33316 14714
rect 33070 14660 33076 14662
rect 33132 14660 33156 14662
rect 33212 14660 33236 14662
rect 33292 14660 33316 14662
rect 33372 14660 33378 14662
rect 33070 14651 33378 14660
rect 3010 14172 3318 14181
rect 3010 14170 3016 14172
rect 3072 14170 3096 14172
rect 3152 14170 3176 14172
rect 3232 14170 3256 14172
rect 3312 14170 3318 14172
rect 3072 14118 3074 14170
rect 3254 14118 3256 14170
rect 3010 14116 3016 14118
rect 3072 14116 3096 14118
rect 3152 14116 3176 14118
rect 3232 14116 3256 14118
rect 3312 14116 3318 14118
rect 3010 14107 3318 14116
rect 33730 14172 34038 14181
rect 33730 14170 33736 14172
rect 33792 14170 33816 14172
rect 33872 14170 33896 14172
rect 33952 14170 33976 14172
rect 34032 14170 34038 14172
rect 33792 14118 33794 14170
rect 33974 14118 33976 14170
rect 33730 14116 33736 14118
rect 33792 14116 33816 14118
rect 33872 14116 33896 14118
rect 33952 14116 33976 14118
rect 34032 14116 34038 14118
rect 33730 14107 34038 14116
rect 2350 13628 2658 13637
rect 2350 13626 2356 13628
rect 2412 13626 2436 13628
rect 2492 13626 2516 13628
rect 2572 13626 2596 13628
rect 2652 13626 2658 13628
rect 2412 13574 2414 13626
rect 2594 13574 2596 13626
rect 2350 13572 2356 13574
rect 2412 13572 2436 13574
rect 2492 13572 2516 13574
rect 2572 13572 2596 13574
rect 2652 13572 2658 13574
rect 2350 13563 2658 13572
rect 33070 13628 33378 13637
rect 33070 13626 33076 13628
rect 33132 13626 33156 13628
rect 33212 13626 33236 13628
rect 33292 13626 33316 13628
rect 33372 13626 33378 13628
rect 33132 13574 33134 13626
rect 33314 13574 33316 13626
rect 33070 13572 33076 13574
rect 33132 13572 33156 13574
rect 33212 13572 33236 13574
rect 33292 13572 33316 13574
rect 33372 13572 33378 13574
rect 33070 13563 33378 13572
rect 3010 13084 3318 13093
rect 3010 13082 3016 13084
rect 3072 13082 3096 13084
rect 3152 13082 3176 13084
rect 3232 13082 3256 13084
rect 3312 13082 3318 13084
rect 3072 13030 3074 13082
rect 3254 13030 3256 13082
rect 3010 13028 3016 13030
rect 3072 13028 3096 13030
rect 3152 13028 3176 13030
rect 3232 13028 3256 13030
rect 3312 13028 3318 13030
rect 3010 13019 3318 13028
rect 33730 13084 34038 13093
rect 33730 13082 33736 13084
rect 33792 13082 33816 13084
rect 33872 13082 33896 13084
rect 33952 13082 33976 13084
rect 34032 13082 34038 13084
rect 33792 13030 33794 13082
rect 33974 13030 33976 13082
rect 33730 13028 33736 13030
rect 33792 13028 33816 13030
rect 33872 13028 33896 13030
rect 33952 13028 33976 13030
rect 34032 13028 34038 13030
rect 33730 13019 34038 13028
rect 2350 12540 2658 12549
rect 2350 12538 2356 12540
rect 2412 12538 2436 12540
rect 2492 12538 2516 12540
rect 2572 12538 2596 12540
rect 2652 12538 2658 12540
rect 2412 12486 2414 12538
rect 2594 12486 2596 12538
rect 2350 12484 2356 12486
rect 2412 12484 2436 12486
rect 2492 12484 2516 12486
rect 2572 12484 2596 12486
rect 2652 12484 2658 12486
rect 2350 12475 2658 12484
rect 33070 12540 33378 12549
rect 33070 12538 33076 12540
rect 33132 12538 33156 12540
rect 33212 12538 33236 12540
rect 33292 12538 33316 12540
rect 33372 12538 33378 12540
rect 33132 12486 33134 12538
rect 33314 12486 33316 12538
rect 33070 12484 33076 12486
rect 33132 12484 33156 12486
rect 33212 12484 33236 12486
rect 33292 12484 33316 12486
rect 33372 12484 33378 12486
rect 33070 12475 33378 12484
rect 3010 11996 3318 12005
rect 3010 11994 3016 11996
rect 3072 11994 3096 11996
rect 3152 11994 3176 11996
rect 3232 11994 3256 11996
rect 3312 11994 3318 11996
rect 3072 11942 3074 11994
rect 3254 11942 3256 11994
rect 3010 11940 3016 11942
rect 3072 11940 3096 11942
rect 3152 11940 3176 11942
rect 3232 11940 3256 11942
rect 3312 11940 3318 11942
rect 3010 11931 3318 11940
rect 33730 11996 34038 12005
rect 33730 11994 33736 11996
rect 33792 11994 33816 11996
rect 33872 11994 33896 11996
rect 33952 11994 33976 11996
rect 34032 11994 34038 11996
rect 33792 11942 33794 11994
rect 33974 11942 33976 11994
rect 33730 11940 33736 11942
rect 33792 11940 33816 11942
rect 33872 11940 33896 11942
rect 33952 11940 33976 11942
rect 34032 11940 34038 11942
rect 33730 11931 34038 11940
rect 2350 11452 2658 11461
rect 2350 11450 2356 11452
rect 2412 11450 2436 11452
rect 2492 11450 2516 11452
rect 2572 11450 2596 11452
rect 2652 11450 2658 11452
rect 2412 11398 2414 11450
rect 2594 11398 2596 11450
rect 2350 11396 2356 11398
rect 2412 11396 2436 11398
rect 2492 11396 2516 11398
rect 2572 11396 2596 11398
rect 2652 11396 2658 11398
rect 2350 11387 2658 11396
rect 33070 11452 33378 11461
rect 33070 11450 33076 11452
rect 33132 11450 33156 11452
rect 33212 11450 33236 11452
rect 33292 11450 33316 11452
rect 33372 11450 33378 11452
rect 33132 11398 33134 11450
rect 33314 11398 33316 11450
rect 33070 11396 33076 11398
rect 33132 11396 33156 11398
rect 33212 11396 33236 11398
rect 33292 11396 33316 11398
rect 33372 11396 33378 11398
rect 33070 11387 33378 11396
rect 3010 10908 3318 10917
rect 3010 10906 3016 10908
rect 3072 10906 3096 10908
rect 3152 10906 3176 10908
rect 3232 10906 3256 10908
rect 3312 10906 3318 10908
rect 3072 10854 3074 10906
rect 3254 10854 3256 10906
rect 3010 10852 3016 10854
rect 3072 10852 3096 10854
rect 3152 10852 3176 10854
rect 3232 10852 3256 10854
rect 3312 10852 3318 10854
rect 3010 10843 3318 10852
rect 33730 10908 34038 10917
rect 33730 10906 33736 10908
rect 33792 10906 33816 10908
rect 33872 10906 33896 10908
rect 33952 10906 33976 10908
rect 34032 10906 34038 10908
rect 33792 10854 33794 10906
rect 33974 10854 33976 10906
rect 33730 10852 33736 10854
rect 33792 10852 33816 10854
rect 33872 10852 33896 10854
rect 33952 10852 33976 10854
rect 34032 10852 34038 10854
rect 33730 10843 34038 10852
rect 2350 10364 2658 10373
rect 2350 10362 2356 10364
rect 2412 10362 2436 10364
rect 2492 10362 2516 10364
rect 2572 10362 2596 10364
rect 2652 10362 2658 10364
rect 2412 10310 2414 10362
rect 2594 10310 2596 10362
rect 2350 10308 2356 10310
rect 2412 10308 2436 10310
rect 2492 10308 2516 10310
rect 2572 10308 2596 10310
rect 2652 10308 2658 10310
rect 2350 10299 2658 10308
rect 33070 10364 33378 10373
rect 33070 10362 33076 10364
rect 33132 10362 33156 10364
rect 33212 10362 33236 10364
rect 33292 10362 33316 10364
rect 33372 10362 33378 10364
rect 33132 10310 33134 10362
rect 33314 10310 33316 10362
rect 33070 10308 33076 10310
rect 33132 10308 33156 10310
rect 33212 10308 33236 10310
rect 33292 10308 33316 10310
rect 33372 10308 33378 10310
rect 33070 10299 33378 10308
rect 3010 9820 3318 9829
rect 3010 9818 3016 9820
rect 3072 9818 3096 9820
rect 3152 9818 3176 9820
rect 3232 9818 3256 9820
rect 3312 9818 3318 9820
rect 3072 9766 3074 9818
rect 3254 9766 3256 9818
rect 3010 9764 3016 9766
rect 3072 9764 3096 9766
rect 3152 9764 3176 9766
rect 3232 9764 3256 9766
rect 3312 9764 3318 9766
rect 3010 9755 3318 9764
rect 33730 9820 34038 9829
rect 33730 9818 33736 9820
rect 33792 9818 33816 9820
rect 33872 9818 33896 9820
rect 33952 9818 33976 9820
rect 34032 9818 34038 9820
rect 33792 9766 33794 9818
rect 33974 9766 33976 9818
rect 33730 9764 33736 9766
rect 33792 9764 33816 9766
rect 33872 9764 33896 9766
rect 33952 9764 33976 9766
rect 34032 9764 34038 9766
rect 33730 9755 34038 9764
rect 2350 9276 2658 9285
rect 2350 9274 2356 9276
rect 2412 9274 2436 9276
rect 2492 9274 2516 9276
rect 2572 9274 2596 9276
rect 2652 9274 2658 9276
rect 2412 9222 2414 9274
rect 2594 9222 2596 9274
rect 2350 9220 2356 9222
rect 2412 9220 2436 9222
rect 2492 9220 2516 9222
rect 2572 9220 2596 9222
rect 2652 9220 2658 9222
rect 2350 9211 2658 9220
rect 33070 9276 33378 9285
rect 33070 9274 33076 9276
rect 33132 9274 33156 9276
rect 33212 9274 33236 9276
rect 33292 9274 33316 9276
rect 33372 9274 33378 9276
rect 33132 9222 33134 9274
rect 33314 9222 33316 9274
rect 33070 9220 33076 9222
rect 33132 9220 33156 9222
rect 33212 9220 33236 9222
rect 33292 9220 33316 9222
rect 33372 9220 33378 9222
rect 33070 9211 33378 9220
rect 3010 8732 3318 8741
rect 3010 8730 3016 8732
rect 3072 8730 3096 8732
rect 3152 8730 3176 8732
rect 3232 8730 3256 8732
rect 3312 8730 3318 8732
rect 3072 8678 3074 8730
rect 3254 8678 3256 8730
rect 3010 8676 3016 8678
rect 3072 8676 3096 8678
rect 3152 8676 3176 8678
rect 3232 8676 3256 8678
rect 3312 8676 3318 8678
rect 3010 8667 3318 8676
rect 33730 8732 34038 8741
rect 33730 8730 33736 8732
rect 33792 8730 33816 8732
rect 33872 8730 33896 8732
rect 33952 8730 33976 8732
rect 34032 8730 34038 8732
rect 33792 8678 33794 8730
rect 33974 8678 33976 8730
rect 33730 8676 33736 8678
rect 33792 8676 33816 8678
rect 33872 8676 33896 8678
rect 33952 8676 33976 8678
rect 34032 8676 34038 8678
rect 33730 8667 34038 8676
rect 2350 8188 2658 8197
rect 2350 8186 2356 8188
rect 2412 8186 2436 8188
rect 2492 8186 2516 8188
rect 2572 8186 2596 8188
rect 2652 8186 2658 8188
rect 2412 8134 2414 8186
rect 2594 8134 2596 8186
rect 2350 8132 2356 8134
rect 2412 8132 2436 8134
rect 2492 8132 2516 8134
rect 2572 8132 2596 8134
rect 2652 8132 2658 8134
rect 2350 8123 2658 8132
rect 33070 8188 33378 8197
rect 33070 8186 33076 8188
rect 33132 8186 33156 8188
rect 33212 8186 33236 8188
rect 33292 8186 33316 8188
rect 33372 8186 33378 8188
rect 33132 8134 33134 8186
rect 33314 8134 33316 8186
rect 33070 8132 33076 8134
rect 33132 8132 33156 8134
rect 33212 8132 33236 8134
rect 33292 8132 33316 8134
rect 33372 8132 33378 8134
rect 33070 8123 33378 8132
rect 3010 7644 3318 7653
rect 3010 7642 3016 7644
rect 3072 7642 3096 7644
rect 3152 7642 3176 7644
rect 3232 7642 3256 7644
rect 3312 7642 3318 7644
rect 3072 7590 3074 7642
rect 3254 7590 3256 7642
rect 3010 7588 3016 7590
rect 3072 7588 3096 7590
rect 3152 7588 3176 7590
rect 3232 7588 3256 7590
rect 3312 7588 3318 7590
rect 3010 7579 3318 7588
rect 33730 7644 34038 7653
rect 33730 7642 33736 7644
rect 33792 7642 33816 7644
rect 33872 7642 33896 7644
rect 33952 7642 33976 7644
rect 34032 7642 34038 7644
rect 33792 7590 33794 7642
rect 33974 7590 33976 7642
rect 33730 7588 33736 7590
rect 33792 7588 33816 7590
rect 33872 7588 33896 7590
rect 33952 7588 33976 7590
rect 34032 7588 34038 7590
rect 33730 7579 34038 7588
rect 2350 7100 2658 7109
rect 2350 7098 2356 7100
rect 2412 7098 2436 7100
rect 2492 7098 2516 7100
rect 2572 7098 2596 7100
rect 2652 7098 2658 7100
rect 2412 7046 2414 7098
rect 2594 7046 2596 7098
rect 2350 7044 2356 7046
rect 2412 7044 2436 7046
rect 2492 7044 2516 7046
rect 2572 7044 2596 7046
rect 2652 7044 2658 7046
rect 2350 7035 2658 7044
rect 33070 7100 33378 7109
rect 33070 7098 33076 7100
rect 33132 7098 33156 7100
rect 33212 7098 33236 7100
rect 33292 7098 33316 7100
rect 33372 7098 33378 7100
rect 33132 7046 33134 7098
rect 33314 7046 33316 7098
rect 33070 7044 33076 7046
rect 33132 7044 33156 7046
rect 33212 7044 33236 7046
rect 33292 7044 33316 7046
rect 33372 7044 33378 7046
rect 33070 7035 33378 7044
rect 3010 6556 3318 6565
rect 3010 6554 3016 6556
rect 3072 6554 3096 6556
rect 3152 6554 3176 6556
rect 3232 6554 3256 6556
rect 3312 6554 3318 6556
rect 3072 6502 3074 6554
rect 3254 6502 3256 6554
rect 3010 6500 3016 6502
rect 3072 6500 3096 6502
rect 3152 6500 3176 6502
rect 3232 6500 3256 6502
rect 3312 6500 3318 6502
rect 3010 6491 3318 6500
rect 33730 6556 34038 6565
rect 33730 6554 33736 6556
rect 33792 6554 33816 6556
rect 33872 6554 33896 6556
rect 33952 6554 33976 6556
rect 34032 6554 34038 6556
rect 33792 6502 33794 6554
rect 33974 6502 33976 6554
rect 33730 6500 33736 6502
rect 33792 6500 33816 6502
rect 33872 6500 33896 6502
rect 33952 6500 33976 6502
rect 34032 6500 34038 6502
rect 33730 6491 34038 6500
rect 2350 6012 2658 6021
rect 2350 6010 2356 6012
rect 2412 6010 2436 6012
rect 2492 6010 2516 6012
rect 2572 6010 2596 6012
rect 2652 6010 2658 6012
rect 2412 5958 2414 6010
rect 2594 5958 2596 6010
rect 2350 5956 2356 5958
rect 2412 5956 2436 5958
rect 2492 5956 2516 5958
rect 2572 5956 2596 5958
rect 2652 5956 2658 5958
rect 2350 5947 2658 5956
rect 33070 6012 33378 6021
rect 33070 6010 33076 6012
rect 33132 6010 33156 6012
rect 33212 6010 33236 6012
rect 33292 6010 33316 6012
rect 33372 6010 33378 6012
rect 33132 5958 33134 6010
rect 33314 5958 33316 6010
rect 33070 5956 33076 5958
rect 33132 5956 33156 5958
rect 33212 5956 33236 5958
rect 33292 5956 33316 5958
rect 33372 5956 33378 5958
rect 33070 5947 33378 5956
rect 3010 5468 3318 5477
rect 3010 5466 3016 5468
rect 3072 5466 3096 5468
rect 3152 5466 3176 5468
rect 3232 5466 3256 5468
rect 3312 5466 3318 5468
rect 3072 5414 3074 5466
rect 3254 5414 3256 5466
rect 3010 5412 3016 5414
rect 3072 5412 3096 5414
rect 3152 5412 3176 5414
rect 3232 5412 3256 5414
rect 3312 5412 3318 5414
rect 3010 5403 3318 5412
rect 33730 5468 34038 5477
rect 33730 5466 33736 5468
rect 33792 5466 33816 5468
rect 33872 5466 33896 5468
rect 33952 5466 33976 5468
rect 34032 5466 34038 5468
rect 33792 5414 33794 5466
rect 33974 5414 33976 5466
rect 33730 5412 33736 5414
rect 33792 5412 33816 5414
rect 33872 5412 33896 5414
rect 33952 5412 33976 5414
rect 34032 5412 34038 5414
rect 33730 5403 34038 5412
rect 2350 4924 2658 4933
rect 2350 4922 2356 4924
rect 2412 4922 2436 4924
rect 2492 4922 2516 4924
rect 2572 4922 2596 4924
rect 2652 4922 2658 4924
rect 2412 4870 2414 4922
rect 2594 4870 2596 4922
rect 2350 4868 2356 4870
rect 2412 4868 2436 4870
rect 2492 4868 2516 4870
rect 2572 4868 2596 4870
rect 2652 4868 2658 4870
rect 2350 4859 2658 4868
rect 33070 4924 33378 4933
rect 33070 4922 33076 4924
rect 33132 4922 33156 4924
rect 33212 4922 33236 4924
rect 33292 4922 33316 4924
rect 33372 4922 33378 4924
rect 33132 4870 33134 4922
rect 33314 4870 33316 4922
rect 33070 4868 33076 4870
rect 33132 4868 33156 4870
rect 33212 4868 33236 4870
rect 33292 4868 33316 4870
rect 33372 4868 33378 4870
rect 33070 4859 33378 4868
rect 3010 4380 3318 4389
rect 3010 4378 3016 4380
rect 3072 4378 3096 4380
rect 3152 4378 3176 4380
rect 3232 4378 3256 4380
rect 3312 4378 3318 4380
rect 3072 4326 3074 4378
rect 3254 4326 3256 4378
rect 3010 4324 3016 4326
rect 3072 4324 3096 4326
rect 3152 4324 3176 4326
rect 3232 4324 3256 4326
rect 3312 4324 3318 4326
rect 3010 4315 3318 4324
rect 33730 4380 34038 4389
rect 33730 4378 33736 4380
rect 33792 4378 33816 4380
rect 33872 4378 33896 4380
rect 33952 4378 33976 4380
rect 34032 4378 34038 4380
rect 33792 4326 33794 4378
rect 33974 4326 33976 4378
rect 33730 4324 33736 4326
rect 33792 4324 33816 4326
rect 33872 4324 33896 4326
rect 33952 4324 33976 4326
rect 34032 4324 34038 4326
rect 33730 4315 34038 4324
rect 2350 3836 2658 3845
rect 2350 3834 2356 3836
rect 2412 3834 2436 3836
rect 2492 3834 2516 3836
rect 2572 3834 2596 3836
rect 2652 3834 2658 3836
rect 2412 3782 2414 3834
rect 2594 3782 2596 3834
rect 2350 3780 2356 3782
rect 2412 3780 2436 3782
rect 2492 3780 2516 3782
rect 2572 3780 2596 3782
rect 2652 3780 2658 3782
rect 2350 3771 2658 3780
rect 33070 3836 33378 3845
rect 33070 3834 33076 3836
rect 33132 3834 33156 3836
rect 33212 3834 33236 3836
rect 33292 3834 33316 3836
rect 33372 3834 33378 3836
rect 33132 3782 33134 3834
rect 33314 3782 33316 3834
rect 33070 3780 33076 3782
rect 33132 3780 33156 3782
rect 33212 3780 33236 3782
rect 33292 3780 33316 3782
rect 33372 3780 33378 3782
rect 33070 3771 33378 3780
rect 3010 3292 3318 3301
rect 3010 3290 3016 3292
rect 3072 3290 3096 3292
rect 3152 3290 3176 3292
rect 3232 3290 3256 3292
rect 3312 3290 3318 3292
rect 3072 3238 3074 3290
rect 3254 3238 3256 3290
rect 3010 3236 3016 3238
rect 3072 3236 3096 3238
rect 3152 3236 3176 3238
rect 3232 3236 3256 3238
rect 3312 3236 3318 3238
rect 3010 3227 3318 3236
rect 33730 3292 34038 3301
rect 33730 3290 33736 3292
rect 33792 3290 33816 3292
rect 33872 3290 33896 3292
rect 33952 3290 33976 3292
rect 34032 3290 34038 3292
rect 33792 3238 33794 3290
rect 33974 3238 33976 3290
rect 33730 3236 33736 3238
rect 33792 3236 33816 3238
rect 33872 3236 33896 3238
rect 33952 3236 33976 3238
rect 34032 3236 34038 3238
rect 33730 3227 34038 3236
rect 2350 2748 2658 2757
rect 2350 2746 2356 2748
rect 2412 2746 2436 2748
rect 2492 2746 2516 2748
rect 2572 2746 2596 2748
rect 2652 2746 2658 2748
rect 2412 2694 2414 2746
rect 2594 2694 2596 2746
rect 2350 2692 2356 2694
rect 2412 2692 2436 2694
rect 2492 2692 2516 2694
rect 2572 2692 2596 2694
rect 2652 2692 2658 2694
rect 2350 2683 2658 2692
rect 33070 2748 33378 2757
rect 33070 2746 33076 2748
rect 33132 2746 33156 2748
rect 33212 2746 33236 2748
rect 33292 2746 33316 2748
rect 33372 2746 33378 2748
rect 33132 2694 33134 2746
rect 33314 2694 33316 2746
rect 33070 2692 33076 2694
rect 33132 2692 33156 2694
rect 33212 2692 33236 2694
rect 33292 2692 33316 2694
rect 33372 2692 33378 2694
rect 33070 2683 33378 2692
rect 3010 2204 3318 2213
rect 3010 2202 3016 2204
rect 3072 2202 3096 2204
rect 3152 2202 3176 2204
rect 3232 2202 3256 2204
rect 3312 2202 3318 2204
rect 3072 2150 3074 2202
rect 3254 2150 3256 2202
rect 3010 2148 3016 2150
rect 3072 2148 3096 2150
rect 3152 2148 3176 2150
rect 3232 2148 3256 2150
rect 3312 2148 3318 2150
rect 3010 2139 3318 2148
rect 33730 2204 34038 2213
rect 33730 2202 33736 2204
rect 33792 2202 33816 2204
rect 33872 2202 33896 2204
rect 33952 2202 33976 2204
rect 34032 2202 34038 2204
rect 33792 2150 33794 2202
rect 33974 2150 33976 2202
rect 33730 2148 33736 2150
rect 33792 2148 33816 2150
rect 33872 2148 33896 2150
rect 33952 2148 33976 2150
rect 34032 2148 34038 2150
rect 33730 2139 34038 2148
<< via2 >>
rect 3016 57690 3072 57692
rect 3096 57690 3152 57692
rect 3176 57690 3232 57692
rect 3256 57690 3312 57692
rect 3016 57638 3062 57690
rect 3062 57638 3072 57690
rect 3096 57638 3126 57690
rect 3126 57638 3138 57690
rect 3138 57638 3152 57690
rect 3176 57638 3190 57690
rect 3190 57638 3202 57690
rect 3202 57638 3232 57690
rect 3256 57638 3266 57690
rect 3266 57638 3312 57690
rect 3016 57636 3072 57638
rect 3096 57636 3152 57638
rect 3176 57636 3232 57638
rect 3256 57636 3312 57638
rect 2356 57146 2412 57148
rect 2436 57146 2492 57148
rect 2516 57146 2572 57148
rect 2596 57146 2652 57148
rect 2356 57094 2402 57146
rect 2402 57094 2412 57146
rect 2436 57094 2466 57146
rect 2466 57094 2478 57146
rect 2478 57094 2492 57146
rect 2516 57094 2530 57146
rect 2530 57094 2542 57146
rect 2542 57094 2572 57146
rect 2596 57094 2606 57146
rect 2606 57094 2652 57146
rect 2356 57092 2412 57094
rect 2436 57092 2492 57094
rect 2516 57092 2572 57094
rect 2596 57092 2652 57094
rect 3016 56602 3072 56604
rect 3096 56602 3152 56604
rect 3176 56602 3232 56604
rect 3256 56602 3312 56604
rect 3016 56550 3062 56602
rect 3062 56550 3072 56602
rect 3096 56550 3126 56602
rect 3126 56550 3138 56602
rect 3138 56550 3152 56602
rect 3176 56550 3190 56602
rect 3190 56550 3202 56602
rect 3202 56550 3232 56602
rect 3256 56550 3266 56602
rect 3266 56550 3312 56602
rect 3016 56548 3072 56550
rect 3096 56548 3152 56550
rect 3176 56548 3232 56550
rect 3256 56548 3312 56550
rect 2356 56058 2412 56060
rect 2436 56058 2492 56060
rect 2516 56058 2572 56060
rect 2596 56058 2652 56060
rect 2356 56006 2402 56058
rect 2402 56006 2412 56058
rect 2436 56006 2466 56058
rect 2466 56006 2478 56058
rect 2478 56006 2492 56058
rect 2516 56006 2530 56058
rect 2530 56006 2542 56058
rect 2542 56006 2572 56058
rect 2596 56006 2606 56058
rect 2606 56006 2652 56058
rect 2356 56004 2412 56006
rect 2436 56004 2492 56006
rect 2516 56004 2572 56006
rect 2596 56004 2652 56006
rect 33736 57690 33792 57692
rect 33816 57690 33872 57692
rect 33896 57690 33952 57692
rect 33976 57690 34032 57692
rect 33736 57638 33782 57690
rect 33782 57638 33792 57690
rect 33816 57638 33846 57690
rect 33846 57638 33858 57690
rect 33858 57638 33872 57690
rect 33896 57638 33910 57690
rect 33910 57638 33922 57690
rect 33922 57638 33952 57690
rect 33976 57638 33986 57690
rect 33986 57638 34032 57690
rect 33736 57636 33792 57638
rect 33816 57636 33872 57638
rect 33896 57636 33952 57638
rect 33976 57636 34032 57638
rect 3016 55514 3072 55516
rect 3096 55514 3152 55516
rect 3176 55514 3232 55516
rect 3256 55514 3312 55516
rect 3016 55462 3062 55514
rect 3062 55462 3072 55514
rect 3096 55462 3126 55514
rect 3126 55462 3138 55514
rect 3138 55462 3152 55514
rect 3176 55462 3190 55514
rect 3190 55462 3202 55514
rect 3202 55462 3232 55514
rect 3256 55462 3266 55514
rect 3266 55462 3312 55514
rect 3016 55460 3072 55462
rect 3096 55460 3152 55462
rect 3176 55460 3232 55462
rect 3256 55460 3312 55462
rect 2356 54970 2412 54972
rect 2436 54970 2492 54972
rect 2516 54970 2572 54972
rect 2596 54970 2652 54972
rect 2356 54918 2402 54970
rect 2402 54918 2412 54970
rect 2436 54918 2466 54970
rect 2466 54918 2478 54970
rect 2478 54918 2492 54970
rect 2516 54918 2530 54970
rect 2530 54918 2542 54970
rect 2542 54918 2572 54970
rect 2596 54918 2606 54970
rect 2606 54918 2652 54970
rect 2356 54916 2412 54918
rect 2436 54916 2492 54918
rect 2516 54916 2572 54918
rect 2596 54916 2652 54918
rect 3016 54426 3072 54428
rect 3096 54426 3152 54428
rect 3176 54426 3232 54428
rect 3256 54426 3312 54428
rect 3016 54374 3062 54426
rect 3062 54374 3072 54426
rect 3096 54374 3126 54426
rect 3126 54374 3138 54426
rect 3138 54374 3152 54426
rect 3176 54374 3190 54426
rect 3190 54374 3202 54426
rect 3202 54374 3232 54426
rect 3256 54374 3266 54426
rect 3266 54374 3312 54426
rect 3016 54372 3072 54374
rect 3096 54372 3152 54374
rect 3176 54372 3232 54374
rect 3256 54372 3312 54374
rect 17406 56480 17462 56536
rect 17222 55564 17224 55584
rect 17224 55564 17276 55584
rect 17276 55564 17278 55584
rect 17222 55528 17278 55564
rect 16946 55256 17002 55312
rect 17314 55256 17370 55312
rect 2356 53882 2412 53884
rect 2436 53882 2492 53884
rect 2516 53882 2572 53884
rect 2596 53882 2652 53884
rect 2356 53830 2402 53882
rect 2402 53830 2412 53882
rect 2436 53830 2466 53882
rect 2466 53830 2478 53882
rect 2478 53830 2492 53882
rect 2516 53830 2530 53882
rect 2530 53830 2542 53882
rect 2542 53830 2572 53882
rect 2596 53830 2606 53882
rect 2606 53830 2652 53882
rect 2356 53828 2412 53830
rect 2436 53828 2492 53830
rect 2516 53828 2572 53830
rect 2596 53828 2652 53830
rect 3016 53338 3072 53340
rect 3096 53338 3152 53340
rect 3176 53338 3232 53340
rect 3256 53338 3312 53340
rect 3016 53286 3062 53338
rect 3062 53286 3072 53338
rect 3096 53286 3126 53338
rect 3126 53286 3138 53338
rect 3138 53286 3152 53338
rect 3176 53286 3190 53338
rect 3190 53286 3202 53338
rect 3202 53286 3232 53338
rect 3256 53286 3266 53338
rect 3266 53286 3312 53338
rect 3016 53284 3072 53286
rect 3096 53284 3152 53286
rect 3176 53284 3232 53286
rect 3256 53284 3312 53286
rect 19890 56480 19946 56536
rect 19614 55528 19670 55584
rect 20534 55820 20590 55856
rect 20534 55800 20536 55820
rect 20536 55800 20588 55820
rect 20588 55800 20590 55820
rect 21914 55836 21916 55856
rect 21916 55836 21968 55856
rect 21968 55836 21970 55856
rect 21914 55800 21970 55836
rect 22834 55528 22890 55584
rect 33076 57146 33132 57148
rect 33156 57146 33212 57148
rect 33236 57146 33292 57148
rect 33316 57146 33372 57148
rect 33076 57094 33122 57146
rect 33122 57094 33132 57146
rect 33156 57094 33186 57146
rect 33186 57094 33198 57146
rect 33198 57094 33212 57146
rect 33236 57094 33250 57146
rect 33250 57094 33262 57146
rect 33262 57094 33292 57146
rect 33316 57094 33326 57146
rect 33326 57094 33372 57146
rect 33076 57092 33132 57094
rect 33156 57092 33212 57094
rect 33236 57092 33292 57094
rect 33316 57092 33372 57094
rect 33736 56602 33792 56604
rect 33816 56602 33872 56604
rect 33896 56602 33952 56604
rect 33976 56602 34032 56604
rect 33736 56550 33782 56602
rect 33782 56550 33792 56602
rect 33816 56550 33846 56602
rect 33846 56550 33858 56602
rect 33858 56550 33872 56602
rect 33896 56550 33910 56602
rect 33910 56550 33922 56602
rect 33922 56550 33952 56602
rect 33976 56550 33986 56602
rect 33986 56550 34032 56602
rect 33736 56548 33792 56550
rect 33816 56548 33872 56550
rect 33896 56548 33952 56550
rect 33976 56548 34032 56550
rect 33076 56058 33132 56060
rect 33156 56058 33212 56060
rect 33236 56058 33292 56060
rect 33316 56058 33372 56060
rect 33076 56006 33122 56058
rect 33122 56006 33132 56058
rect 33156 56006 33186 56058
rect 33186 56006 33198 56058
rect 33198 56006 33212 56058
rect 33236 56006 33250 56058
rect 33250 56006 33262 56058
rect 33262 56006 33292 56058
rect 33316 56006 33326 56058
rect 33326 56006 33372 56058
rect 33076 56004 33132 56006
rect 33156 56004 33212 56006
rect 33236 56004 33292 56006
rect 33316 56004 33372 56006
rect 33736 55514 33792 55516
rect 33816 55514 33872 55516
rect 33896 55514 33952 55516
rect 33976 55514 34032 55516
rect 33736 55462 33782 55514
rect 33782 55462 33792 55514
rect 33816 55462 33846 55514
rect 33846 55462 33858 55514
rect 33858 55462 33872 55514
rect 33896 55462 33910 55514
rect 33910 55462 33922 55514
rect 33922 55462 33952 55514
rect 33976 55462 33986 55514
rect 33986 55462 34032 55514
rect 33736 55460 33792 55462
rect 33816 55460 33872 55462
rect 33896 55460 33952 55462
rect 33976 55460 34032 55462
rect 33076 54970 33132 54972
rect 33156 54970 33212 54972
rect 33236 54970 33292 54972
rect 33316 54970 33372 54972
rect 33076 54918 33122 54970
rect 33122 54918 33132 54970
rect 33156 54918 33186 54970
rect 33186 54918 33198 54970
rect 33198 54918 33212 54970
rect 33236 54918 33250 54970
rect 33250 54918 33262 54970
rect 33262 54918 33292 54970
rect 33316 54918 33326 54970
rect 33326 54918 33372 54970
rect 33076 54916 33132 54918
rect 33156 54916 33212 54918
rect 33236 54916 33292 54918
rect 33316 54916 33372 54918
rect 33736 54426 33792 54428
rect 33816 54426 33872 54428
rect 33896 54426 33952 54428
rect 33976 54426 34032 54428
rect 33736 54374 33782 54426
rect 33782 54374 33792 54426
rect 33816 54374 33846 54426
rect 33846 54374 33858 54426
rect 33858 54374 33872 54426
rect 33896 54374 33910 54426
rect 33910 54374 33922 54426
rect 33922 54374 33952 54426
rect 33976 54374 33986 54426
rect 33986 54374 34032 54426
rect 33736 54372 33792 54374
rect 33816 54372 33872 54374
rect 33896 54372 33952 54374
rect 33976 54372 34032 54374
rect 33076 53882 33132 53884
rect 33156 53882 33212 53884
rect 33236 53882 33292 53884
rect 33316 53882 33372 53884
rect 33076 53830 33122 53882
rect 33122 53830 33132 53882
rect 33156 53830 33186 53882
rect 33186 53830 33198 53882
rect 33198 53830 33212 53882
rect 33236 53830 33250 53882
rect 33250 53830 33262 53882
rect 33262 53830 33292 53882
rect 33316 53830 33326 53882
rect 33326 53830 33372 53882
rect 33076 53828 33132 53830
rect 33156 53828 33212 53830
rect 33236 53828 33292 53830
rect 33316 53828 33372 53830
rect 33736 53338 33792 53340
rect 33816 53338 33872 53340
rect 33896 53338 33952 53340
rect 33976 53338 34032 53340
rect 33736 53286 33782 53338
rect 33782 53286 33792 53338
rect 33816 53286 33846 53338
rect 33846 53286 33858 53338
rect 33858 53286 33872 53338
rect 33896 53286 33910 53338
rect 33910 53286 33922 53338
rect 33922 53286 33952 53338
rect 33976 53286 33986 53338
rect 33986 53286 34032 53338
rect 33736 53284 33792 53286
rect 33816 53284 33872 53286
rect 33896 53284 33952 53286
rect 33976 53284 34032 53286
rect 2356 52794 2412 52796
rect 2436 52794 2492 52796
rect 2516 52794 2572 52796
rect 2596 52794 2652 52796
rect 2356 52742 2402 52794
rect 2402 52742 2412 52794
rect 2436 52742 2466 52794
rect 2466 52742 2478 52794
rect 2478 52742 2492 52794
rect 2516 52742 2530 52794
rect 2530 52742 2542 52794
rect 2542 52742 2572 52794
rect 2596 52742 2606 52794
rect 2606 52742 2652 52794
rect 2356 52740 2412 52742
rect 2436 52740 2492 52742
rect 2516 52740 2572 52742
rect 2596 52740 2652 52742
rect 33076 52794 33132 52796
rect 33156 52794 33212 52796
rect 33236 52794 33292 52796
rect 33316 52794 33372 52796
rect 33076 52742 33122 52794
rect 33122 52742 33132 52794
rect 33156 52742 33186 52794
rect 33186 52742 33198 52794
rect 33198 52742 33212 52794
rect 33236 52742 33250 52794
rect 33250 52742 33262 52794
rect 33262 52742 33292 52794
rect 33316 52742 33326 52794
rect 33326 52742 33372 52794
rect 33076 52740 33132 52742
rect 33156 52740 33212 52742
rect 33236 52740 33292 52742
rect 33316 52740 33372 52742
rect 3016 52250 3072 52252
rect 3096 52250 3152 52252
rect 3176 52250 3232 52252
rect 3256 52250 3312 52252
rect 3016 52198 3062 52250
rect 3062 52198 3072 52250
rect 3096 52198 3126 52250
rect 3126 52198 3138 52250
rect 3138 52198 3152 52250
rect 3176 52198 3190 52250
rect 3190 52198 3202 52250
rect 3202 52198 3232 52250
rect 3256 52198 3266 52250
rect 3266 52198 3312 52250
rect 3016 52196 3072 52198
rect 3096 52196 3152 52198
rect 3176 52196 3232 52198
rect 3256 52196 3312 52198
rect 33736 52250 33792 52252
rect 33816 52250 33872 52252
rect 33896 52250 33952 52252
rect 33976 52250 34032 52252
rect 33736 52198 33782 52250
rect 33782 52198 33792 52250
rect 33816 52198 33846 52250
rect 33846 52198 33858 52250
rect 33858 52198 33872 52250
rect 33896 52198 33910 52250
rect 33910 52198 33922 52250
rect 33922 52198 33952 52250
rect 33976 52198 33986 52250
rect 33986 52198 34032 52250
rect 33736 52196 33792 52198
rect 33816 52196 33872 52198
rect 33896 52196 33952 52198
rect 33976 52196 34032 52198
rect 2356 51706 2412 51708
rect 2436 51706 2492 51708
rect 2516 51706 2572 51708
rect 2596 51706 2652 51708
rect 2356 51654 2402 51706
rect 2402 51654 2412 51706
rect 2436 51654 2466 51706
rect 2466 51654 2478 51706
rect 2478 51654 2492 51706
rect 2516 51654 2530 51706
rect 2530 51654 2542 51706
rect 2542 51654 2572 51706
rect 2596 51654 2606 51706
rect 2606 51654 2652 51706
rect 2356 51652 2412 51654
rect 2436 51652 2492 51654
rect 2516 51652 2572 51654
rect 2596 51652 2652 51654
rect 33076 51706 33132 51708
rect 33156 51706 33212 51708
rect 33236 51706 33292 51708
rect 33316 51706 33372 51708
rect 33076 51654 33122 51706
rect 33122 51654 33132 51706
rect 33156 51654 33186 51706
rect 33186 51654 33198 51706
rect 33198 51654 33212 51706
rect 33236 51654 33250 51706
rect 33250 51654 33262 51706
rect 33262 51654 33292 51706
rect 33316 51654 33326 51706
rect 33326 51654 33372 51706
rect 33076 51652 33132 51654
rect 33156 51652 33212 51654
rect 33236 51652 33292 51654
rect 33316 51652 33372 51654
rect 3016 51162 3072 51164
rect 3096 51162 3152 51164
rect 3176 51162 3232 51164
rect 3256 51162 3312 51164
rect 3016 51110 3062 51162
rect 3062 51110 3072 51162
rect 3096 51110 3126 51162
rect 3126 51110 3138 51162
rect 3138 51110 3152 51162
rect 3176 51110 3190 51162
rect 3190 51110 3202 51162
rect 3202 51110 3232 51162
rect 3256 51110 3266 51162
rect 3266 51110 3312 51162
rect 3016 51108 3072 51110
rect 3096 51108 3152 51110
rect 3176 51108 3232 51110
rect 3256 51108 3312 51110
rect 33736 51162 33792 51164
rect 33816 51162 33872 51164
rect 33896 51162 33952 51164
rect 33976 51162 34032 51164
rect 33736 51110 33782 51162
rect 33782 51110 33792 51162
rect 33816 51110 33846 51162
rect 33846 51110 33858 51162
rect 33858 51110 33872 51162
rect 33896 51110 33910 51162
rect 33910 51110 33922 51162
rect 33922 51110 33952 51162
rect 33976 51110 33986 51162
rect 33986 51110 34032 51162
rect 33736 51108 33792 51110
rect 33816 51108 33872 51110
rect 33896 51108 33952 51110
rect 33976 51108 34032 51110
rect 2356 50618 2412 50620
rect 2436 50618 2492 50620
rect 2516 50618 2572 50620
rect 2596 50618 2652 50620
rect 2356 50566 2402 50618
rect 2402 50566 2412 50618
rect 2436 50566 2466 50618
rect 2466 50566 2478 50618
rect 2478 50566 2492 50618
rect 2516 50566 2530 50618
rect 2530 50566 2542 50618
rect 2542 50566 2572 50618
rect 2596 50566 2606 50618
rect 2606 50566 2652 50618
rect 2356 50564 2412 50566
rect 2436 50564 2492 50566
rect 2516 50564 2572 50566
rect 2596 50564 2652 50566
rect 33076 50618 33132 50620
rect 33156 50618 33212 50620
rect 33236 50618 33292 50620
rect 33316 50618 33372 50620
rect 33076 50566 33122 50618
rect 33122 50566 33132 50618
rect 33156 50566 33186 50618
rect 33186 50566 33198 50618
rect 33198 50566 33212 50618
rect 33236 50566 33250 50618
rect 33250 50566 33262 50618
rect 33262 50566 33292 50618
rect 33316 50566 33326 50618
rect 33326 50566 33372 50618
rect 33076 50564 33132 50566
rect 33156 50564 33212 50566
rect 33236 50564 33292 50566
rect 33316 50564 33372 50566
rect 3016 50074 3072 50076
rect 3096 50074 3152 50076
rect 3176 50074 3232 50076
rect 3256 50074 3312 50076
rect 3016 50022 3062 50074
rect 3062 50022 3072 50074
rect 3096 50022 3126 50074
rect 3126 50022 3138 50074
rect 3138 50022 3152 50074
rect 3176 50022 3190 50074
rect 3190 50022 3202 50074
rect 3202 50022 3232 50074
rect 3256 50022 3266 50074
rect 3266 50022 3312 50074
rect 3016 50020 3072 50022
rect 3096 50020 3152 50022
rect 3176 50020 3232 50022
rect 3256 50020 3312 50022
rect 33736 50074 33792 50076
rect 33816 50074 33872 50076
rect 33896 50074 33952 50076
rect 33976 50074 34032 50076
rect 33736 50022 33782 50074
rect 33782 50022 33792 50074
rect 33816 50022 33846 50074
rect 33846 50022 33858 50074
rect 33858 50022 33872 50074
rect 33896 50022 33910 50074
rect 33910 50022 33922 50074
rect 33922 50022 33952 50074
rect 33976 50022 33986 50074
rect 33986 50022 34032 50074
rect 33736 50020 33792 50022
rect 33816 50020 33872 50022
rect 33896 50020 33952 50022
rect 33976 50020 34032 50022
rect 2356 49530 2412 49532
rect 2436 49530 2492 49532
rect 2516 49530 2572 49532
rect 2596 49530 2652 49532
rect 2356 49478 2402 49530
rect 2402 49478 2412 49530
rect 2436 49478 2466 49530
rect 2466 49478 2478 49530
rect 2478 49478 2492 49530
rect 2516 49478 2530 49530
rect 2530 49478 2542 49530
rect 2542 49478 2572 49530
rect 2596 49478 2606 49530
rect 2606 49478 2652 49530
rect 2356 49476 2412 49478
rect 2436 49476 2492 49478
rect 2516 49476 2572 49478
rect 2596 49476 2652 49478
rect 33076 49530 33132 49532
rect 33156 49530 33212 49532
rect 33236 49530 33292 49532
rect 33316 49530 33372 49532
rect 33076 49478 33122 49530
rect 33122 49478 33132 49530
rect 33156 49478 33186 49530
rect 33186 49478 33198 49530
rect 33198 49478 33212 49530
rect 33236 49478 33250 49530
rect 33250 49478 33262 49530
rect 33262 49478 33292 49530
rect 33316 49478 33326 49530
rect 33326 49478 33372 49530
rect 33076 49476 33132 49478
rect 33156 49476 33212 49478
rect 33236 49476 33292 49478
rect 33316 49476 33372 49478
rect 3016 48986 3072 48988
rect 3096 48986 3152 48988
rect 3176 48986 3232 48988
rect 3256 48986 3312 48988
rect 3016 48934 3062 48986
rect 3062 48934 3072 48986
rect 3096 48934 3126 48986
rect 3126 48934 3138 48986
rect 3138 48934 3152 48986
rect 3176 48934 3190 48986
rect 3190 48934 3202 48986
rect 3202 48934 3232 48986
rect 3256 48934 3266 48986
rect 3266 48934 3312 48986
rect 3016 48932 3072 48934
rect 3096 48932 3152 48934
rect 3176 48932 3232 48934
rect 3256 48932 3312 48934
rect 33736 48986 33792 48988
rect 33816 48986 33872 48988
rect 33896 48986 33952 48988
rect 33976 48986 34032 48988
rect 33736 48934 33782 48986
rect 33782 48934 33792 48986
rect 33816 48934 33846 48986
rect 33846 48934 33858 48986
rect 33858 48934 33872 48986
rect 33896 48934 33910 48986
rect 33910 48934 33922 48986
rect 33922 48934 33952 48986
rect 33976 48934 33986 48986
rect 33986 48934 34032 48986
rect 33736 48932 33792 48934
rect 33816 48932 33872 48934
rect 33896 48932 33952 48934
rect 33976 48932 34032 48934
rect 2356 48442 2412 48444
rect 2436 48442 2492 48444
rect 2516 48442 2572 48444
rect 2596 48442 2652 48444
rect 2356 48390 2402 48442
rect 2402 48390 2412 48442
rect 2436 48390 2466 48442
rect 2466 48390 2478 48442
rect 2478 48390 2492 48442
rect 2516 48390 2530 48442
rect 2530 48390 2542 48442
rect 2542 48390 2572 48442
rect 2596 48390 2606 48442
rect 2606 48390 2652 48442
rect 2356 48388 2412 48390
rect 2436 48388 2492 48390
rect 2516 48388 2572 48390
rect 2596 48388 2652 48390
rect 33076 48442 33132 48444
rect 33156 48442 33212 48444
rect 33236 48442 33292 48444
rect 33316 48442 33372 48444
rect 33076 48390 33122 48442
rect 33122 48390 33132 48442
rect 33156 48390 33186 48442
rect 33186 48390 33198 48442
rect 33198 48390 33212 48442
rect 33236 48390 33250 48442
rect 33250 48390 33262 48442
rect 33262 48390 33292 48442
rect 33316 48390 33326 48442
rect 33326 48390 33372 48442
rect 33076 48388 33132 48390
rect 33156 48388 33212 48390
rect 33236 48388 33292 48390
rect 33316 48388 33372 48390
rect 3016 47898 3072 47900
rect 3096 47898 3152 47900
rect 3176 47898 3232 47900
rect 3256 47898 3312 47900
rect 3016 47846 3062 47898
rect 3062 47846 3072 47898
rect 3096 47846 3126 47898
rect 3126 47846 3138 47898
rect 3138 47846 3152 47898
rect 3176 47846 3190 47898
rect 3190 47846 3202 47898
rect 3202 47846 3232 47898
rect 3256 47846 3266 47898
rect 3266 47846 3312 47898
rect 3016 47844 3072 47846
rect 3096 47844 3152 47846
rect 3176 47844 3232 47846
rect 3256 47844 3312 47846
rect 33736 47898 33792 47900
rect 33816 47898 33872 47900
rect 33896 47898 33952 47900
rect 33976 47898 34032 47900
rect 33736 47846 33782 47898
rect 33782 47846 33792 47898
rect 33816 47846 33846 47898
rect 33846 47846 33858 47898
rect 33858 47846 33872 47898
rect 33896 47846 33910 47898
rect 33910 47846 33922 47898
rect 33922 47846 33952 47898
rect 33976 47846 33986 47898
rect 33986 47846 34032 47898
rect 33736 47844 33792 47846
rect 33816 47844 33872 47846
rect 33896 47844 33952 47846
rect 33976 47844 34032 47846
rect 2356 47354 2412 47356
rect 2436 47354 2492 47356
rect 2516 47354 2572 47356
rect 2596 47354 2652 47356
rect 2356 47302 2402 47354
rect 2402 47302 2412 47354
rect 2436 47302 2466 47354
rect 2466 47302 2478 47354
rect 2478 47302 2492 47354
rect 2516 47302 2530 47354
rect 2530 47302 2542 47354
rect 2542 47302 2572 47354
rect 2596 47302 2606 47354
rect 2606 47302 2652 47354
rect 2356 47300 2412 47302
rect 2436 47300 2492 47302
rect 2516 47300 2572 47302
rect 2596 47300 2652 47302
rect 33076 47354 33132 47356
rect 33156 47354 33212 47356
rect 33236 47354 33292 47356
rect 33316 47354 33372 47356
rect 33076 47302 33122 47354
rect 33122 47302 33132 47354
rect 33156 47302 33186 47354
rect 33186 47302 33198 47354
rect 33198 47302 33212 47354
rect 33236 47302 33250 47354
rect 33250 47302 33262 47354
rect 33262 47302 33292 47354
rect 33316 47302 33326 47354
rect 33326 47302 33372 47354
rect 33076 47300 33132 47302
rect 33156 47300 33212 47302
rect 33236 47300 33292 47302
rect 33316 47300 33372 47302
rect 3016 46810 3072 46812
rect 3096 46810 3152 46812
rect 3176 46810 3232 46812
rect 3256 46810 3312 46812
rect 3016 46758 3062 46810
rect 3062 46758 3072 46810
rect 3096 46758 3126 46810
rect 3126 46758 3138 46810
rect 3138 46758 3152 46810
rect 3176 46758 3190 46810
rect 3190 46758 3202 46810
rect 3202 46758 3232 46810
rect 3256 46758 3266 46810
rect 3266 46758 3312 46810
rect 3016 46756 3072 46758
rect 3096 46756 3152 46758
rect 3176 46756 3232 46758
rect 3256 46756 3312 46758
rect 33736 46810 33792 46812
rect 33816 46810 33872 46812
rect 33896 46810 33952 46812
rect 33976 46810 34032 46812
rect 33736 46758 33782 46810
rect 33782 46758 33792 46810
rect 33816 46758 33846 46810
rect 33846 46758 33858 46810
rect 33858 46758 33872 46810
rect 33896 46758 33910 46810
rect 33910 46758 33922 46810
rect 33922 46758 33952 46810
rect 33976 46758 33986 46810
rect 33986 46758 34032 46810
rect 33736 46756 33792 46758
rect 33816 46756 33872 46758
rect 33896 46756 33952 46758
rect 33976 46756 34032 46758
rect 2356 46266 2412 46268
rect 2436 46266 2492 46268
rect 2516 46266 2572 46268
rect 2596 46266 2652 46268
rect 2356 46214 2402 46266
rect 2402 46214 2412 46266
rect 2436 46214 2466 46266
rect 2466 46214 2478 46266
rect 2478 46214 2492 46266
rect 2516 46214 2530 46266
rect 2530 46214 2542 46266
rect 2542 46214 2572 46266
rect 2596 46214 2606 46266
rect 2606 46214 2652 46266
rect 2356 46212 2412 46214
rect 2436 46212 2492 46214
rect 2516 46212 2572 46214
rect 2596 46212 2652 46214
rect 33076 46266 33132 46268
rect 33156 46266 33212 46268
rect 33236 46266 33292 46268
rect 33316 46266 33372 46268
rect 33076 46214 33122 46266
rect 33122 46214 33132 46266
rect 33156 46214 33186 46266
rect 33186 46214 33198 46266
rect 33198 46214 33212 46266
rect 33236 46214 33250 46266
rect 33250 46214 33262 46266
rect 33262 46214 33292 46266
rect 33316 46214 33326 46266
rect 33326 46214 33372 46266
rect 33076 46212 33132 46214
rect 33156 46212 33212 46214
rect 33236 46212 33292 46214
rect 33316 46212 33372 46214
rect 3016 45722 3072 45724
rect 3096 45722 3152 45724
rect 3176 45722 3232 45724
rect 3256 45722 3312 45724
rect 3016 45670 3062 45722
rect 3062 45670 3072 45722
rect 3096 45670 3126 45722
rect 3126 45670 3138 45722
rect 3138 45670 3152 45722
rect 3176 45670 3190 45722
rect 3190 45670 3202 45722
rect 3202 45670 3232 45722
rect 3256 45670 3266 45722
rect 3266 45670 3312 45722
rect 3016 45668 3072 45670
rect 3096 45668 3152 45670
rect 3176 45668 3232 45670
rect 3256 45668 3312 45670
rect 33736 45722 33792 45724
rect 33816 45722 33872 45724
rect 33896 45722 33952 45724
rect 33976 45722 34032 45724
rect 33736 45670 33782 45722
rect 33782 45670 33792 45722
rect 33816 45670 33846 45722
rect 33846 45670 33858 45722
rect 33858 45670 33872 45722
rect 33896 45670 33910 45722
rect 33910 45670 33922 45722
rect 33922 45670 33952 45722
rect 33976 45670 33986 45722
rect 33986 45670 34032 45722
rect 33736 45668 33792 45670
rect 33816 45668 33872 45670
rect 33896 45668 33952 45670
rect 33976 45668 34032 45670
rect 49054 55256 49110 55312
rect 2356 45178 2412 45180
rect 2436 45178 2492 45180
rect 2516 45178 2572 45180
rect 2596 45178 2652 45180
rect 2356 45126 2402 45178
rect 2402 45126 2412 45178
rect 2436 45126 2466 45178
rect 2466 45126 2478 45178
rect 2478 45126 2492 45178
rect 2516 45126 2530 45178
rect 2530 45126 2542 45178
rect 2542 45126 2572 45178
rect 2596 45126 2606 45178
rect 2606 45126 2652 45178
rect 2356 45124 2412 45126
rect 2436 45124 2492 45126
rect 2516 45124 2572 45126
rect 2596 45124 2652 45126
rect 33076 45178 33132 45180
rect 33156 45178 33212 45180
rect 33236 45178 33292 45180
rect 33316 45178 33372 45180
rect 33076 45126 33122 45178
rect 33122 45126 33132 45178
rect 33156 45126 33186 45178
rect 33186 45126 33198 45178
rect 33198 45126 33212 45178
rect 33236 45126 33250 45178
rect 33250 45126 33262 45178
rect 33262 45126 33292 45178
rect 33316 45126 33326 45178
rect 33326 45126 33372 45178
rect 33076 45124 33132 45126
rect 33156 45124 33212 45126
rect 33236 45124 33292 45126
rect 33316 45124 33372 45126
rect 3016 44634 3072 44636
rect 3096 44634 3152 44636
rect 3176 44634 3232 44636
rect 3256 44634 3312 44636
rect 3016 44582 3062 44634
rect 3062 44582 3072 44634
rect 3096 44582 3126 44634
rect 3126 44582 3138 44634
rect 3138 44582 3152 44634
rect 3176 44582 3190 44634
rect 3190 44582 3202 44634
rect 3202 44582 3232 44634
rect 3256 44582 3266 44634
rect 3266 44582 3312 44634
rect 3016 44580 3072 44582
rect 3096 44580 3152 44582
rect 3176 44580 3232 44582
rect 3256 44580 3312 44582
rect 33736 44634 33792 44636
rect 33816 44634 33872 44636
rect 33896 44634 33952 44636
rect 33976 44634 34032 44636
rect 33736 44582 33782 44634
rect 33782 44582 33792 44634
rect 33816 44582 33846 44634
rect 33846 44582 33858 44634
rect 33858 44582 33872 44634
rect 33896 44582 33910 44634
rect 33910 44582 33922 44634
rect 33922 44582 33952 44634
rect 33976 44582 33986 44634
rect 33986 44582 34032 44634
rect 33736 44580 33792 44582
rect 33816 44580 33872 44582
rect 33896 44580 33952 44582
rect 33976 44580 34032 44582
rect 2356 44090 2412 44092
rect 2436 44090 2492 44092
rect 2516 44090 2572 44092
rect 2596 44090 2652 44092
rect 2356 44038 2402 44090
rect 2402 44038 2412 44090
rect 2436 44038 2466 44090
rect 2466 44038 2478 44090
rect 2478 44038 2492 44090
rect 2516 44038 2530 44090
rect 2530 44038 2542 44090
rect 2542 44038 2572 44090
rect 2596 44038 2606 44090
rect 2606 44038 2652 44090
rect 2356 44036 2412 44038
rect 2436 44036 2492 44038
rect 2516 44036 2572 44038
rect 2596 44036 2652 44038
rect 33076 44090 33132 44092
rect 33156 44090 33212 44092
rect 33236 44090 33292 44092
rect 33316 44090 33372 44092
rect 33076 44038 33122 44090
rect 33122 44038 33132 44090
rect 33156 44038 33186 44090
rect 33186 44038 33198 44090
rect 33198 44038 33212 44090
rect 33236 44038 33250 44090
rect 33250 44038 33262 44090
rect 33262 44038 33292 44090
rect 33316 44038 33326 44090
rect 33326 44038 33372 44090
rect 33076 44036 33132 44038
rect 33156 44036 33212 44038
rect 33236 44036 33292 44038
rect 33316 44036 33372 44038
rect 3016 43546 3072 43548
rect 3096 43546 3152 43548
rect 3176 43546 3232 43548
rect 3256 43546 3312 43548
rect 3016 43494 3062 43546
rect 3062 43494 3072 43546
rect 3096 43494 3126 43546
rect 3126 43494 3138 43546
rect 3138 43494 3152 43546
rect 3176 43494 3190 43546
rect 3190 43494 3202 43546
rect 3202 43494 3232 43546
rect 3256 43494 3266 43546
rect 3266 43494 3312 43546
rect 3016 43492 3072 43494
rect 3096 43492 3152 43494
rect 3176 43492 3232 43494
rect 3256 43492 3312 43494
rect 33736 43546 33792 43548
rect 33816 43546 33872 43548
rect 33896 43546 33952 43548
rect 33976 43546 34032 43548
rect 33736 43494 33782 43546
rect 33782 43494 33792 43546
rect 33816 43494 33846 43546
rect 33846 43494 33858 43546
rect 33858 43494 33872 43546
rect 33896 43494 33910 43546
rect 33910 43494 33922 43546
rect 33922 43494 33952 43546
rect 33976 43494 33986 43546
rect 33986 43494 34032 43546
rect 33736 43492 33792 43494
rect 33816 43492 33872 43494
rect 33896 43492 33952 43494
rect 33976 43492 34032 43494
rect 2356 43002 2412 43004
rect 2436 43002 2492 43004
rect 2516 43002 2572 43004
rect 2596 43002 2652 43004
rect 2356 42950 2402 43002
rect 2402 42950 2412 43002
rect 2436 42950 2466 43002
rect 2466 42950 2478 43002
rect 2478 42950 2492 43002
rect 2516 42950 2530 43002
rect 2530 42950 2542 43002
rect 2542 42950 2572 43002
rect 2596 42950 2606 43002
rect 2606 42950 2652 43002
rect 2356 42948 2412 42950
rect 2436 42948 2492 42950
rect 2516 42948 2572 42950
rect 2596 42948 2652 42950
rect 33076 43002 33132 43004
rect 33156 43002 33212 43004
rect 33236 43002 33292 43004
rect 33316 43002 33372 43004
rect 33076 42950 33122 43002
rect 33122 42950 33132 43002
rect 33156 42950 33186 43002
rect 33186 42950 33198 43002
rect 33198 42950 33212 43002
rect 33236 42950 33250 43002
rect 33250 42950 33262 43002
rect 33262 42950 33292 43002
rect 33316 42950 33326 43002
rect 33326 42950 33372 43002
rect 33076 42948 33132 42950
rect 33156 42948 33212 42950
rect 33236 42948 33292 42950
rect 33316 42948 33372 42950
rect 3016 42458 3072 42460
rect 3096 42458 3152 42460
rect 3176 42458 3232 42460
rect 3256 42458 3312 42460
rect 3016 42406 3062 42458
rect 3062 42406 3072 42458
rect 3096 42406 3126 42458
rect 3126 42406 3138 42458
rect 3138 42406 3152 42458
rect 3176 42406 3190 42458
rect 3190 42406 3202 42458
rect 3202 42406 3232 42458
rect 3256 42406 3266 42458
rect 3266 42406 3312 42458
rect 3016 42404 3072 42406
rect 3096 42404 3152 42406
rect 3176 42404 3232 42406
rect 3256 42404 3312 42406
rect 33736 42458 33792 42460
rect 33816 42458 33872 42460
rect 33896 42458 33952 42460
rect 33976 42458 34032 42460
rect 33736 42406 33782 42458
rect 33782 42406 33792 42458
rect 33816 42406 33846 42458
rect 33846 42406 33858 42458
rect 33858 42406 33872 42458
rect 33896 42406 33910 42458
rect 33910 42406 33922 42458
rect 33922 42406 33952 42458
rect 33976 42406 33986 42458
rect 33986 42406 34032 42458
rect 33736 42404 33792 42406
rect 33816 42404 33872 42406
rect 33896 42404 33952 42406
rect 33976 42404 34032 42406
rect 2356 41914 2412 41916
rect 2436 41914 2492 41916
rect 2516 41914 2572 41916
rect 2596 41914 2652 41916
rect 2356 41862 2402 41914
rect 2402 41862 2412 41914
rect 2436 41862 2466 41914
rect 2466 41862 2478 41914
rect 2478 41862 2492 41914
rect 2516 41862 2530 41914
rect 2530 41862 2542 41914
rect 2542 41862 2572 41914
rect 2596 41862 2606 41914
rect 2606 41862 2652 41914
rect 2356 41860 2412 41862
rect 2436 41860 2492 41862
rect 2516 41860 2572 41862
rect 2596 41860 2652 41862
rect 33076 41914 33132 41916
rect 33156 41914 33212 41916
rect 33236 41914 33292 41916
rect 33316 41914 33372 41916
rect 33076 41862 33122 41914
rect 33122 41862 33132 41914
rect 33156 41862 33186 41914
rect 33186 41862 33198 41914
rect 33198 41862 33212 41914
rect 33236 41862 33250 41914
rect 33250 41862 33262 41914
rect 33262 41862 33292 41914
rect 33316 41862 33326 41914
rect 33326 41862 33372 41914
rect 33076 41860 33132 41862
rect 33156 41860 33212 41862
rect 33236 41860 33292 41862
rect 33316 41860 33372 41862
rect 3016 41370 3072 41372
rect 3096 41370 3152 41372
rect 3176 41370 3232 41372
rect 3256 41370 3312 41372
rect 3016 41318 3062 41370
rect 3062 41318 3072 41370
rect 3096 41318 3126 41370
rect 3126 41318 3138 41370
rect 3138 41318 3152 41370
rect 3176 41318 3190 41370
rect 3190 41318 3202 41370
rect 3202 41318 3232 41370
rect 3256 41318 3266 41370
rect 3266 41318 3312 41370
rect 3016 41316 3072 41318
rect 3096 41316 3152 41318
rect 3176 41316 3232 41318
rect 3256 41316 3312 41318
rect 33736 41370 33792 41372
rect 33816 41370 33872 41372
rect 33896 41370 33952 41372
rect 33976 41370 34032 41372
rect 33736 41318 33782 41370
rect 33782 41318 33792 41370
rect 33816 41318 33846 41370
rect 33846 41318 33858 41370
rect 33858 41318 33872 41370
rect 33896 41318 33910 41370
rect 33910 41318 33922 41370
rect 33922 41318 33952 41370
rect 33976 41318 33986 41370
rect 33986 41318 34032 41370
rect 33736 41316 33792 41318
rect 33816 41316 33872 41318
rect 33896 41316 33952 41318
rect 33976 41316 34032 41318
rect 2356 40826 2412 40828
rect 2436 40826 2492 40828
rect 2516 40826 2572 40828
rect 2596 40826 2652 40828
rect 2356 40774 2402 40826
rect 2402 40774 2412 40826
rect 2436 40774 2466 40826
rect 2466 40774 2478 40826
rect 2478 40774 2492 40826
rect 2516 40774 2530 40826
rect 2530 40774 2542 40826
rect 2542 40774 2572 40826
rect 2596 40774 2606 40826
rect 2606 40774 2652 40826
rect 2356 40772 2412 40774
rect 2436 40772 2492 40774
rect 2516 40772 2572 40774
rect 2596 40772 2652 40774
rect 33076 40826 33132 40828
rect 33156 40826 33212 40828
rect 33236 40826 33292 40828
rect 33316 40826 33372 40828
rect 33076 40774 33122 40826
rect 33122 40774 33132 40826
rect 33156 40774 33186 40826
rect 33186 40774 33198 40826
rect 33198 40774 33212 40826
rect 33236 40774 33250 40826
rect 33250 40774 33262 40826
rect 33262 40774 33292 40826
rect 33316 40774 33326 40826
rect 33326 40774 33372 40826
rect 33076 40772 33132 40774
rect 33156 40772 33212 40774
rect 33236 40772 33292 40774
rect 33316 40772 33372 40774
rect 3016 40282 3072 40284
rect 3096 40282 3152 40284
rect 3176 40282 3232 40284
rect 3256 40282 3312 40284
rect 3016 40230 3062 40282
rect 3062 40230 3072 40282
rect 3096 40230 3126 40282
rect 3126 40230 3138 40282
rect 3138 40230 3152 40282
rect 3176 40230 3190 40282
rect 3190 40230 3202 40282
rect 3202 40230 3232 40282
rect 3256 40230 3266 40282
rect 3266 40230 3312 40282
rect 3016 40228 3072 40230
rect 3096 40228 3152 40230
rect 3176 40228 3232 40230
rect 3256 40228 3312 40230
rect 33736 40282 33792 40284
rect 33816 40282 33872 40284
rect 33896 40282 33952 40284
rect 33976 40282 34032 40284
rect 33736 40230 33782 40282
rect 33782 40230 33792 40282
rect 33816 40230 33846 40282
rect 33846 40230 33858 40282
rect 33858 40230 33872 40282
rect 33896 40230 33910 40282
rect 33910 40230 33922 40282
rect 33922 40230 33952 40282
rect 33976 40230 33986 40282
rect 33986 40230 34032 40282
rect 33736 40228 33792 40230
rect 33816 40228 33872 40230
rect 33896 40228 33952 40230
rect 33976 40228 34032 40230
rect 2356 39738 2412 39740
rect 2436 39738 2492 39740
rect 2516 39738 2572 39740
rect 2596 39738 2652 39740
rect 2356 39686 2402 39738
rect 2402 39686 2412 39738
rect 2436 39686 2466 39738
rect 2466 39686 2478 39738
rect 2478 39686 2492 39738
rect 2516 39686 2530 39738
rect 2530 39686 2542 39738
rect 2542 39686 2572 39738
rect 2596 39686 2606 39738
rect 2606 39686 2652 39738
rect 2356 39684 2412 39686
rect 2436 39684 2492 39686
rect 2516 39684 2572 39686
rect 2596 39684 2652 39686
rect 33076 39738 33132 39740
rect 33156 39738 33212 39740
rect 33236 39738 33292 39740
rect 33316 39738 33372 39740
rect 33076 39686 33122 39738
rect 33122 39686 33132 39738
rect 33156 39686 33186 39738
rect 33186 39686 33198 39738
rect 33198 39686 33212 39738
rect 33236 39686 33250 39738
rect 33250 39686 33262 39738
rect 33262 39686 33292 39738
rect 33316 39686 33326 39738
rect 33326 39686 33372 39738
rect 33076 39684 33132 39686
rect 33156 39684 33212 39686
rect 33236 39684 33292 39686
rect 33316 39684 33372 39686
rect 3016 39194 3072 39196
rect 3096 39194 3152 39196
rect 3176 39194 3232 39196
rect 3256 39194 3312 39196
rect 3016 39142 3062 39194
rect 3062 39142 3072 39194
rect 3096 39142 3126 39194
rect 3126 39142 3138 39194
rect 3138 39142 3152 39194
rect 3176 39142 3190 39194
rect 3190 39142 3202 39194
rect 3202 39142 3232 39194
rect 3256 39142 3266 39194
rect 3266 39142 3312 39194
rect 3016 39140 3072 39142
rect 3096 39140 3152 39142
rect 3176 39140 3232 39142
rect 3256 39140 3312 39142
rect 33736 39194 33792 39196
rect 33816 39194 33872 39196
rect 33896 39194 33952 39196
rect 33976 39194 34032 39196
rect 33736 39142 33782 39194
rect 33782 39142 33792 39194
rect 33816 39142 33846 39194
rect 33846 39142 33858 39194
rect 33858 39142 33872 39194
rect 33896 39142 33910 39194
rect 33910 39142 33922 39194
rect 33922 39142 33952 39194
rect 33976 39142 33986 39194
rect 33986 39142 34032 39194
rect 33736 39140 33792 39142
rect 33816 39140 33872 39142
rect 33896 39140 33952 39142
rect 33976 39140 34032 39142
rect 2356 38650 2412 38652
rect 2436 38650 2492 38652
rect 2516 38650 2572 38652
rect 2596 38650 2652 38652
rect 2356 38598 2402 38650
rect 2402 38598 2412 38650
rect 2436 38598 2466 38650
rect 2466 38598 2478 38650
rect 2478 38598 2492 38650
rect 2516 38598 2530 38650
rect 2530 38598 2542 38650
rect 2542 38598 2572 38650
rect 2596 38598 2606 38650
rect 2606 38598 2652 38650
rect 2356 38596 2412 38598
rect 2436 38596 2492 38598
rect 2516 38596 2572 38598
rect 2596 38596 2652 38598
rect 33076 38650 33132 38652
rect 33156 38650 33212 38652
rect 33236 38650 33292 38652
rect 33316 38650 33372 38652
rect 33076 38598 33122 38650
rect 33122 38598 33132 38650
rect 33156 38598 33186 38650
rect 33186 38598 33198 38650
rect 33198 38598 33212 38650
rect 33236 38598 33250 38650
rect 33250 38598 33262 38650
rect 33262 38598 33292 38650
rect 33316 38598 33326 38650
rect 33326 38598 33372 38650
rect 33076 38596 33132 38598
rect 33156 38596 33212 38598
rect 33236 38596 33292 38598
rect 33316 38596 33372 38598
rect 3016 38106 3072 38108
rect 3096 38106 3152 38108
rect 3176 38106 3232 38108
rect 3256 38106 3312 38108
rect 3016 38054 3062 38106
rect 3062 38054 3072 38106
rect 3096 38054 3126 38106
rect 3126 38054 3138 38106
rect 3138 38054 3152 38106
rect 3176 38054 3190 38106
rect 3190 38054 3202 38106
rect 3202 38054 3232 38106
rect 3256 38054 3266 38106
rect 3266 38054 3312 38106
rect 3016 38052 3072 38054
rect 3096 38052 3152 38054
rect 3176 38052 3232 38054
rect 3256 38052 3312 38054
rect 33736 38106 33792 38108
rect 33816 38106 33872 38108
rect 33896 38106 33952 38108
rect 33976 38106 34032 38108
rect 33736 38054 33782 38106
rect 33782 38054 33792 38106
rect 33816 38054 33846 38106
rect 33846 38054 33858 38106
rect 33858 38054 33872 38106
rect 33896 38054 33910 38106
rect 33910 38054 33922 38106
rect 33922 38054 33952 38106
rect 33976 38054 33986 38106
rect 33986 38054 34032 38106
rect 33736 38052 33792 38054
rect 33816 38052 33872 38054
rect 33896 38052 33952 38054
rect 33976 38052 34032 38054
rect 2356 37562 2412 37564
rect 2436 37562 2492 37564
rect 2516 37562 2572 37564
rect 2596 37562 2652 37564
rect 2356 37510 2402 37562
rect 2402 37510 2412 37562
rect 2436 37510 2466 37562
rect 2466 37510 2478 37562
rect 2478 37510 2492 37562
rect 2516 37510 2530 37562
rect 2530 37510 2542 37562
rect 2542 37510 2572 37562
rect 2596 37510 2606 37562
rect 2606 37510 2652 37562
rect 2356 37508 2412 37510
rect 2436 37508 2492 37510
rect 2516 37508 2572 37510
rect 2596 37508 2652 37510
rect 33076 37562 33132 37564
rect 33156 37562 33212 37564
rect 33236 37562 33292 37564
rect 33316 37562 33372 37564
rect 33076 37510 33122 37562
rect 33122 37510 33132 37562
rect 33156 37510 33186 37562
rect 33186 37510 33198 37562
rect 33198 37510 33212 37562
rect 33236 37510 33250 37562
rect 33250 37510 33262 37562
rect 33262 37510 33292 37562
rect 33316 37510 33326 37562
rect 33326 37510 33372 37562
rect 33076 37508 33132 37510
rect 33156 37508 33212 37510
rect 33236 37508 33292 37510
rect 33316 37508 33372 37510
rect 3016 37018 3072 37020
rect 3096 37018 3152 37020
rect 3176 37018 3232 37020
rect 3256 37018 3312 37020
rect 3016 36966 3062 37018
rect 3062 36966 3072 37018
rect 3096 36966 3126 37018
rect 3126 36966 3138 37018
rect 3138 36966 3152 37018
rect 3176 36966 3190 37018
rect 3190 36966 3202 37018
rect 3202 36966 3232 37018
rect 3256 36966 3266 37018
rect 3266 36966 3312 37018
rect 3016 36964 3072 36966
rect 3096 36964 3152 36966
rect 3176 36964 3232 36966
rect 3256 36964 3312 36966
rect 33736 37018 33792 37020
rect 33816 37018 33872 37020
rect 33896 37018 33952 37020
rect 33976 37018 34032 37020
rect 33736 36966 33782 37018
rect 33782 36966 33792 37018
rect 33816 36966 33846 37018
rect 33846 36966 33858 37018
rect 33858 36966 33872 37018
rect 33896 36966 33910 37018
rect 33910 36966 33922 37018
rect 33922 36966 33952 37018
rect 33976 36966 33986 37018
rect 33986 36966 34032 37018
rect 33736 36964 33792 36966
rect 33816 36964 33872 36966
rect 33896 36964 33952 36966
rect 33976 36964 34032 36966
rect 2356 36474 2412 36476
rect 2436 36474 2492 36476
rect 2516 36474 2572 36476
rect 2596 36474 2652 36476
rect 2356 36422 2402 36474
rect 2402 36422 2412 36474
rect 2436 36422 2466 36474
rect 2466 36422 2478 36474
rect 2478 36422 2492 36474
rect 2516 36422 2530 36474
rect 2530 36422 2542 36474
rect 2542 36422 2572 36474
rect 2596 36422 2606 36474
rect 2606 36422 2652 36474
rect 2356 36420 2412 36422
rect 2436 36420 2492 36422
rect 2516 36420 2572 36422
rect 2596 36420 2652 36422
rect 33076 36474 33132 36476
rect 33156 36474 33212 36476
rect 33236 36474 33292 36476
rect 33316 36474 33372 36476
rect 33076 36422 33122 36474
rect 33122 36422 33132 36474
rect 33156 36422 33186 36474
rect 33186 36422 33198 36474
rect 33198 36422 33212 36474
rect 33236 36422 33250 36474
rect 33250 36422 33262 36474
rect 33262 36422 33292 36474
rect 33316 36422 33326 36474
rect 33326 36422 33372 36474
rect 33076 36420 33132 36422
rect 33156 36420 33212 36422
rect 33236 36420 33292 36422
rect 33316 36420 33372 36422
rect 3016 35930 3072 35932
rect 3096 35930 3152 35932
rect 3176 35930 3232 35932
rect 3256 35930 3312 35932
rect 3016 35878 3062 35930
rect 3062 35878 3072 35930
rect 3096 35878 3126 35930
rect 3126 35878 3138 35930
rect 3138 35878 3152 35930
rect 3176 35878 3190 35930
rect 3190 35878 3202 35930
rect 3202 35878 3232 35930
rect 3256 35878 3266 35930
rect 3266 35878 3312 35930
rect 3016 35876 3072 35878
rect 3096 35876 3152 35878
rect 3176 35876 3232 35878
rect 3256 35876 3312 35878
rect 33736 35930 33792 35932
rect 33816 35930 33872 35932
rect 33896 35930 33952 35932
rect 33976 35930 34032 35932
rect 33736 35878 33782 35930
rect 33782 35878 33792 35930
rect 33816 35878 33846 35930
rect 33846 35878 33858 35930
rect 33858 35878 33872 35930
rect 33896 35878 33910 35930
rect 33910 35878 33922 35930
rect 33922 35878 33952 35930
rect 33976 35878 33986 35930
rect 33986 35878 34032 35930
rect 33736 35876 33792 35878
rect 33816 35876 33872 35878
rect 33896 35876 33952 35878
rect 33976 35876 34032 35878
rect 2356 35386 2412 35388
rect 2436 35386 2492 35388
rect 2516 35386 2572 35388
rect 2596 35386 2652 35388
rect 2356 35334 2402 35386
rect 2402 35334 2412 35386
rect 2436 35334 2466 35386
rect 2466 35334 2478 35386
rect 2478 35334 2492 35386
rect 2516 35334 2530 35386
rect 2530 35334 2542 35386
rect 2542 35334 2572 35386
rect 2596 35334 2606 35386
rect 2606 35334 2652 35386
rect 2356 35332 2412 35334
rect 2436 35332 2492 35334
rect 2516 35332 2572 35334
rect 2596 35332 2652 35334
rect 33076 35386 33132 35388
rect 33156 35386 33212 35388
rect 33236 35386 33292 35388
rect 33316 35386 33372 35388
rect 33076 35334 33122 35386
rect 33122 35334 33132 35386
rect 33156 35334 33186 35386
rect 33186 35334 33198 35386
rect 33198 35334 33212 35386
rect 33236 35334 33250 35386
rect 33250 35334 33262 35386
rect 33262 35334 33292 35386
rect 33316 35334 33326 35386
rect 33326 35334 33372 35386
rect 33076 35332 33132 35334
rect 33156 35332 33212 35334
rect 33236 35332 33292 35334
rect 33316 35332 33372 35334
rect 3016 34842 3072 34844
rect 3096 34842 3152 34844
rect 3176 34842 3232 34844
rect 3256 34842 3312 34844
rect 3016 34790 3062 34842
rect 3062 34790 3072 34842
rect 3096 34790 3126 34842
rect 3126 34790 3138 34842
rect 3138 34790 3152 34842
rect 3176 34790 3190 34842
rect 3190 34790 3202 34842
rect 3202 34790 3232 34842
rect 3256 34790 3266 34842
rect 3266 34790 3312 34842
rect 3016 34788 3072 34790
rect 3096 34788 3152 34790
rect 3176 34788 3232 34790
rect 3256 34788 3312 34790
rect 33736 34842 33792 34844
rect 33816 34842 33872 34844
rect 33896 34842 33952 34844
rect 33976 34842 34032 34844
rect 33736 34790 33782 34842
rect 33782 34790 33792 34842
rect 33816 34790 33846 34842
rect 33846 34790 33858 34842
rect 33858 34790 33872 34842
rect 33896 34790 33910 34842
rect 33910 34790 33922 34842
rect 33922 34790 33952 34842
rect 33976 34790 33986 34842
rect 33986 34790 34032 34842
rect 33736 34788 33792 34790
rect 33816 34788 33872 34790
rect 33896 34788 33952 34790
rect 33976 34788 34032 34790
rect 2356 34298 2412 34300
rect 2436 34298 2492 34300
rect 2516 34298 2572 34300
rect 2596 34298 2652 34300
rect 2356 34246 2402 34298
rect 2402 34246 2412 34298
rect 2436 34246 2466 34298
rect 2466 34246 2478 34298
rect 2478 34246 2492 34298
rect 2516 34246 2530 34298
rect 2530 34246 2542 34298
rect 2542 34246 2572 34298
rect 2596 34246 2606 34298
rect 2606 34246 2652 34298
rect 2356 34244 2412 34246
rect 2436 34244 2492 34246
rect 2516 34244 2572 34246
rect 2596 34244 2652 34246
rect 33076 34298 33132 34300
rect 33156 34298 33212 34300
rect 33236 34298 33292 34300
rect 33316 34298 33372 34300
rect 33076 34246 33122 34298
rect 33122 34246 33132 34298
rect 33156 34246 33186 34298
rect 33186 34246 33198 34298
rect 33198 34246 33212 34298
rect 33236 34246 33250 34298
rect 33250 34246 33262 34298
rect 33262 34246 33292 34298
rect 33316 34246 33326 34298
rect 33326 34246 33372 34298
rect 33076 34244 33132 34246
rect 33156 34244 33212 34246
rect 33236 34244 33292 34246
rect 33316 34244 33372 34246
rect 3016 33754 3072 33756
rect 3096 33754 3152 33756
rect 3176 33754 3232 33756
rect 3256 33754 3312 33756
rect 3016 33702 3062 33754
rect 3062 33702 3072 33754
rect 3096 33702 3126 33754
rect 3126 33702 3138 33754
rect 3138 33702 3152 33754
rect 3176 33702 3190 33754
rect 3190 33702 3202 33754
rect 3202 33702 3232 33754
rect 3256 33702 3266 33754
rect 3266 33702 3312 33754
rect 3016 33700 3072 33702
rect 3096 33700 3152 33702
rect 3176 33700 3232 33702
rect 3256 33700 3312 33702
rect 33736 33754 33792 33756
rect 33816 33754 33872 33756
rect 33896 33754 33952 33756
rect 33976 33754 34032 33756
rect 33736 33702 33782 33754
rect 33782 33702 33792 33754
rect 33816 33702 33846 33754
rect 33846 33702 33858 33754
rect 33858 33702 33872 33754
rect 33896 33702 33910 33754
rect 33910 33702 33922 33754
rect 33922 33702 33952 33754
rect 33976 33702 33986 33754
rect 33986 33702 34032 33754
rect 33736 33700 33792 33702
rect 33816 33700 33872 33702
rect 33896 33700 33952 33702
rect 33976 33700 34032 33702
rect 2356 33210 2412 33212
rect 2436 33210 2492 33212
rect 2516 33210 2572 33212
rect 2596 33210 2652 33212
rect 2356 33158 2402 33210
rect 2402 33158 2412 33210
rect 2436 33158 2466 33210
rect 2466 33158 2478 33210
rect 2478 33158 2492 33210
rect 2516 33158 2530 33210
rect 2530 33158 2542 33210
rect 2542 33158 2572 33210
rect 2596 33158 2606 33210
rect 2606 33158 2652 33210
rect 2356 33156 2412 33158
rect 2436 33156 2492 33158
rect 2516 33156 2572 33158
rect 2596 33156 2652 33158
rect 33076 33210 33132 33212
rect 33156 33210 33212 33212
rect 33236 33210 33292 33212
rect 33316 33210 33372 33212
rect 33076 33158 33122 33210
rect 33122 33158 33132 33210
rect 33156 33158 33186 33210
rect 33186 33158 33198 33210
rect 33198 33158 33212 33210
rect 33236 33158 33250 33210
rect 33250 33158 33262 33210
rect 33262 33158 33292 33210
rect 33316 33158 33326 33210
rect 33326 33158 33372 33210
rect 33076 33156 33132 33158
rect 33156 33156 33212 33158
rect 33236 33156 33292 33158
rect 33316 33156 33372 33158
rect 3016 32666 3072 32668
rect 3096 32666 3152 32668
rect 3176 32666 3232 32668
rect 3256 32666 3312 32668
rect 3016 32614 3062 32666
rect 3062 32614 3072 32666
rect 3096 32614 3126 32666
rect 3126 32614 3138 32666
rect 3138 32614 3152 32666
rect 3176 32614 3190 32666
rect 3190 32614 3202 32666
rect 3202 32614 3232 32666
rect 3256 32614 3266 32666
rect 3266 32614 3312 32666
rect 3016 32612 3072 32614
rect 3096 32612 3152 32614
rect 3176 32612 3232 32614
rect 3256 32612 3312 32614
rect 33736 32666 33792 32668
rect 33816 32666 33872 32668
rect 33896 32666 33952 32668
rect 33976 32666 34032 32668
rect 33736 32614 33782 32666
rect 33782 32614 33792 32666
rect 33816 32614 33846 32666
rect 33846 32614 33858 32666
rect 33858 32614 33872 32666
rect 33896 32614 33910 32666
rect 33910 32614 33922 32666
rect 33922 32614 33952 32666
rect 33976 32614 33986 32666
rect 33986 32614 34032 32666
rect 33736 32612 33792 32614
rect 33816 32612 33872 32614
rect 33896 32612 33952 32614
rect 33976 32612 34032 32614
rect 2356 32122 2412 32124
rect 2436 32122 2492 32124
rect 2516 32122 2572 32124
rect 2596 32122 2652 32124
rect 2356 32070 2402 32122
rect 2402 32070 2412 32122
rect 2436 32070 2466 32122
rect 2466 32070 2478 32122
rect 2478 32070 2492 32122
rect 2516 32070 2530 32122
rect 2530 32070 2542 32122
rect 2542 32070 2572 32122
rect 2596 32070 2606 32122
rect 2606 32070 2652 32122
rect 2356 32068 2412 32070
rect 2436 32068 2492 32070
rect 2516 32068 2572 32070
rect 2596 32068 2652 32070
rect 33076 32122 33132 32124
rect 33156 32122 33212 32124
rect 33236 32122 33292 32124
rect 33316 32122 33372 32124
rect 33076 32070 33122 32122
rect 33122 32070 33132 32122
rect 33156 32070 33186 32122
rect 33186 32070 33198 32122
rect 33198 32070 33212 32122
rect 33236 32070 33250 32122
rect 33250 32070 33262 32122
rect 33262 32070 33292 32122
rect 33316 32070 33326 32122
rect 33326 32070 33372 32122
rect 33076 32068 33132 32070
rect 33156 32068 33212 32070
rect 33236 32068 33292 32070
rect 33316 32068 33372 32070
rect 3016 31578 3072 31580
rect 3096 31578 3152 31580
rect 3176 31578 3232 31580
rect 3256 31578 3312 31580
rect 3016 31526 3062 31578
rect 3062 31526 3072 31578
rect 3096 31526 3126 31578
rect 3126 31526 3138 31578
rect 3138 31526 3152 31578
rect 3176 31526 3190 31578
rect 3190 31526 3202 31578
rect 3202 31526 3232 31578
rect 3256 31526 3266 31578
rect 3266 31526 3312 31578
rect 3016 31524 3072 31526
rect 3096 31524 3152 31526
rect 3176 31524 3232 31526
rect 3256 31524 3312 31526
rect 33736 31578 33792 31580
rect 33816 31578 33872 31580
rect 33896 31578 33952 31580
rect 33976 31578 34032 31580
rect 33736 31526 33782 31578
rect 33782 31526 33792 31578
rect 33816 31526 33846 31578
rect 33846 31526 33858 31578
rect 33858 31526 33872 31578
rect 33896 31526 33910 31578
rect 33910 31526 33922 31578
rect 33922 31526 33952 31578
rect 33976 31526 33986 31578
rect 33986 31526 34032 31578
rect 33736 31524 33792 31526
rect 33816 31524 33872 31526
rect 33896 31524 33952 31526
rect 33976 31524 34032 31526
rect 2356 31034 2412 31036
rect 2436 31034 2492 31036
rect 2516 31034 2572 31036
rect 2596 31034 2652 31036
rect 2356 30982 2402 31034
rect 2402 30982 2412 31034
rect 2436 30982 2466 31034
rect 2466 30982 2478 31034
rect 2478 30982 2492 31034
rect 2516 30982 2530 31034
rect 2530 30982 2542 31034
rect 2542 30982 2572 31034
rect 2596 30982 2606 31034
rect 2606 30982 2652 31034
rect 2356 30980 2412 30982
rect 2436 30980 2492 30982
rect 2516 30980 2572 30982
rect 2596 30980 2652 30982
rect 33076 31034 33132 31036
rect 33156 31034 33212 31036
rect 33236 31034 33292 31036
rect 33316 31034 33372 31036
rect 33076 30982 33122 31034
rect 33122 30982 33132 31034
rect 33156 30982 33186 31034
rect 33186 30982 33198 31034
rect 33198 30982 33212 31034
rect 33236 30982 33250 31034
rect 33250 30982 33262 31034
rect 33262 30982 33292 31034
rect 33316 30982 33326 31034
rect 33326 30982 33372 31034
rect 33076 30980 33132 30982
rect 33156 30980 33212 30982
rect 33236 30980 33292 30982
rect 33316 30980 33372 30982
rect 3016 30490 3072 30492
rect 3096 30490 3152 30492
rect 3176 30490 3232 30492
rect 3256 30490 3312 30492
rect 3016 30438 3062 30490
rect 3062 30438 3072 30490
rect 3096 30438 3126 30490
rect 3126 30438 3138 30490
rect 3138 30438 3152 30490
rect 3176 30438 3190 30490
rect 3190 30438 3202 30490
rect 3202 30438 3232 30490
rect 3256 30438 3266 30490
rect 3266 30438 3312 30490
rect 3016 30436 3072 30438
rect 3096 30436 3152 30438
rect 3176 30436 3232 30438
rect 3256 30436 3312 30438
rect 33736 30490 33792 30492
rect 33816 30490 33872 30492
rect 33896 30490 33952 30492
rect 33976 30490 34032 30492
rect 33736 30438 33782 30490
rect 33782 30438 33792 30490
rect 33816 30438 33846 30490
rect 33846 30438 33858 30490
rect 33858 30438 33872 30490
rect 33896 30438 33910 30490
rect 33910 30438 33922 30490
rect 33922 30438 33952 30490
rect 33976 30438 33986 30490
rect 33986 30438 34032 30490
rect 33736 30436 33792 30438
rect 33816 30436 33872 30438
rect 33896 30436 33952 30438
rect 33976 30436 34032 30438
rect 2356 29946 2412 29948
rect 2436 29946 2492 29948
rect 2516 29946 2572 29948
rect 2596 29946 2652 29948
rect 2356 29894 2402 29946
rect 2402 29894 2412 29946
rect 2436 29894 2466 29946
rect 2466 29894 2478 29946
rect 2478 29894 2492 29946
rect 2516 29894 2530 29946
rect 2530 29894 2542 29946
rect 2542 29894 2572 29946
rect 2596 29894 2606 29946
rect 2606 29894 2652 29946
rect 2356 29892 2412 29894
rect 2436 29892 2492 29894
rect 2516 29892 2572 29894
rect 2596 29892 2652 29894
rect 33076 29946 33132 29948
rect 33156 29946 33212 29948
rect 33236 29946 33292 29948
rect 33316 29946 33372 29948
rect 33076 29894 33122 29946
rect 33122 29894 33132 29946
rect 33156 29894 33186 29946
rect 33186 29894 33198 29946
rect 33198 29894 33212 29946
rect 33236 29894 33250 29946
rect 33250 29894 33262 29946
rect 33262 29894 33292 29946
rect 33316 29894 33326 29946
rect 33326 29894 33372 29946
rect 33076 29892 33132 29894
rect 33156 29892 33212 29894
rect 33236 29892 33292 29894
rect 33316 29892 33372 29894
rect 3016 29402 3072 29404
rect 3096 29402 3152 29404
rect 3176 29402 3232 29404
rect 3256 29402 3312 29404
rect 3016 29350 3062 29402
rect 3062 29350 3072 29402
rect 3096 29350 3126 29402
rect 3126 29350 3138 29402
rect 3138 29350 3152 29402
rect 3176 29350 3190 29402
rect 3190 29350 3202 29402
rect 3202 29350 3232 29402
rect 3256 29350 3266 29402
rect 3266 29350 3312 29402
rect 3016 29348 3072 29350
rect 3096 29348 3152 29350
rect 3176 29348 3232 29350
rect 3256 29348 3312 29350
rect 33736 29402 33792 29404
rect 33816 29402 33872 29404
rect 33896 29402 33952 29404
rect 33976 29402 34032 29404
rect 33736 29350 33782 29402
rect 33782 29350 33792 29402
rect 33816 29350 33846 29402
rect 33846 29350 33858 29402
rect 33858 29350 33872 29402
rect 33896 29350 33910 29402
rect 33910 29350 33922 29402
rect 33922 29350 33952 29402
rect 33976 29350 33986 29402
rect 33986 29350 34032 29402
rect 33736 29348 33792 29350
rect 33816 29348 33872 29350
rect 33896 29348 33952 29350
rect 33976 29348 34032 29350
rect 2356 28858 2412 28860
rect 2436 28858 2492 28860
rect 2516 28858 2572 28860
rect 2596 28858 2652 28860
rect 2356 28806 2402 28858
rect 2402 28806 2412 28858
rect 2436 28806 2466 28858
rect 2466 28806 2478 28858
rect 2478 28806 2492 28858
rect 2516 28806 2530 28858
rect 2530 28806 2542 28858
rect 2542 28806 2572 28858
rect 2596 28806 2606 28858
rect 2606 28806 2652 28858
rect 2356 28804 2412 28806
rect 2436 28804 2492 28806
rect 2516 28804 2572 28806
rect 2596 28804 2652 28806
rect 33076 28858 33132 28860
rect 33156 28858 33212 28860
rect 33236 28858 33292 28860
rect 33316 28858 33372 28860
rect 33076 28806 33122 28858
rect 33122 28806 33132 28858
rect 33156 28806 33186 28858
rect 33186 28806 33198 28858
rect 33198 28806 33212 28858
rect 33236 28806 33250 28858
rect 33250 28806 33262 28858
rect 33262 28806 33292 28858
rect 33316 28806 33326 28858
rect 33326 28806 33372 28858
rect 33076 28804 33132 28806
rect 33156 28804 33212 28806
rect 33236 28804 33292 28806
rect 33316 28804 33372 28806
rect 3016 28314 3072 28316
rect 3096 28314 3152 28316
rect 3176 28314 3232 28316
rect 3256 28314 3312 28316
rect 3016 28262 3062 28314
rect 3062 28262 3072 28314
rect 3096 28262 3126 28314
rect 3126 28262 3138 28314
rect 3138 28262 3152 28314
rect 3176 28262 3190 28314
rect 3190 28262 3202 28314
rect 3202 28262 3232 28314
rect 3256 28262 3266 28314
rect 3266 28262 3312 28314
rect 3016 28260 3072 28262
rect 3096 28260 3152 28262
rect 3176 28260 3232 28262
rect 3256 28260 3312 28262
rect 33736 28314 33792 28316
rect 33816 28314 33872 28316
rect 33896 28314 33952 28316
rect 33976 28314 34032 28316
rect 33736 28262 33782 28314
rect 33782 28262 33792 28314
rect 33816 28262 33846 28314
rect 33846 28262 33858 28314
rect 33858 28262 33872 28314
rect 33896 28262 33910 28314
rect 33910 28262 33922 28314
rect 33922 28262 33952 28314
rect 33976 28262 33986 28314
rect 33986 28262 34032 28314
rect 33736 28260 33792 28262
rect 33816 28260 33872 28262
rect 33896 28260 33952 28262
rect 33976 28260 34032 28262
rect 2356 27770 2412 27772
rect 2436 27770 2492 27772
rect 2516 27770 2572 27772
rect 2596 27770 2652 27772
rect 2356 27718 2402 27770
rect 2402 27718 2412 27770
rect 2436 27718 2466 27770
rect 2466 27718 2478 27770
rect 2478 27718 2492 27770
rect 2516 27718 2530 27770
rect 2530 27718 2542 27770
rect 2542 27718 2572 27770
rect 2596 27718 2606 27770
rect 2606 27718 2652 27770
rect 2356 27716 2412 27718
rect 2436 27716 2492 27718
rect 2516 27716 2572 27718
rect 2596 27716 2652 27718
rect 33076 27770 33132 27772
rect 33156 27770 33212 27772
rect 33236 27770 33292 27772
rect 33316 27770 33372 27772
rect 33076 27718 33122 27770
rect 33122 27718 33132 27770
rect 33156 27718 33186 27770
rect 33186 27718 33198 27770
rect 33198 27718 33212 27770
rect 33236 27718 33250 27770
rect 33250 27718 33262 27770
rect 33262 27718 33292 27770
rect 33316 27718 33326 27770
rect 33326 27718 33372 27770
rect 33076 27716 33132 27718
rect 33156 27716 33212 27718
rect 33236 27716 33292 27718
rect 33316 27716 33372 27718
rect 3016 27226 3072 27228
rect 3096 27226 3152 27228
rect 3176 27226 3232 27228
rect 3256 27226 3312 27228
rect 3016 27174 3062 27226
rect 3062 27174 3072 27226
rect 3096 27174 3126 27226
rect 3126 27174 3138 27226
rect 3138 27174 3152 27226
rect 3176 27174 3190 27226
rect 3190 27174 3202 27226
rect 3202 27174 3232 27226
rect 3256 27174 3266 27226
rect 3266 27174 3312 27226
rect 3016 27172 3072 27174
rect 3096 27172 3152 27174
rect 3176 27172 3232 27174
rect 3256 27172 3312 27174
rect 33736 27226 33792 27228
rect 33816 27226 33872 27228
rect 33896 27226 33952 27228
rect 33976 27226 34032 27228
rect 33736 27174 33782 27226
rect 33782 27174 33792 27226
rect 33816 27174 33846 27226
rect 33846 27174 33858 27226
rect 33858 27174 33872 27226
rect 33896 27174 33910 27226
rect 33910 27174 33922 27226
rect 33922 27174 33952 27226
rect 33976 27174 33986 27226
rect 33986 27174 34032 27226
rect 33736 27172 33792 27174
rect 33816 27172 33872 27174
rect 33896 27172 33952 27174
rect 33976 27172 34032 27174
rect 2356 26682 2412 26684
rect 2436 26682 2492 26684
rect 2516 26682 2572 26684
rect 2596 26682 2652 26684
rect 2356 26630 2402 26682
rect 2402 26630 2412 26682
rect 2436 26630 2466 26682
rect 2466 26630 2478 26682
rect 2478 26630 2492 26682
rect 2516 26630 2530 26682
rect 2530 26630 2542 26682
rect 2542 26630 2572 26682
rect 2596 26630 2606 26682
rect 2606 26630 2652 26682
rect 2356 26628 2412 26630
rect 2436 26628 2492 26630
rect 2516 26628 2572 26630
rect 2596 26628 2652 26630
rect 33076 26682 33132 26684
rect 33156 26682 33212 26684
rect 33236 26682 33292 26684
rect 33316 26682 33372 26684
rect 33076 26630 33122 26682
rect 33122 26630 33132 26682
rect 33156 26630 33186 26682
rect 33186 26630 33198 26682
rect 33198 26630 33212 26682
rect 33236 26630 33250 26682
rect 33250 26630 33262 26682
rect 33262 26630 33292 26682
rect 33316 26630 33326 26682
rect 33326 26630 33372 26682
rect 33076 26628 33132 26630
rect 33156 26628 33212 26630
rect 33236 26628 33292 26630
rect 33316 26628 33372 26630
rect 3016 26138 3072 26140
rect 3096 26138 3152 26140
rect 3176 26138 3232 26140
rect 3256 26138 3312 26140
rect 3016 26086 3062 26138
rect 3062 26086 3072 26138
rect 3096 26086 3126 26138
rect 3126 26086 3138 26138
rect 3138 26086 3152 26138
rect 3176 26086 3190 26138
rect 3190 26086 3202 26138
rect 3202 26086 3232 26138
rect 3256 26086 3266 26138
rect 3266 26086 3312 26138
rect 3016 26084 3072 26086
rect 3096 26084 3152 26086
rect 3176 26084 3232 26086
rect 3256 26084 3312 26086
rect 33736 26138 33792 26140
rect 33816 26138 33872 26140
rect 33896 26138 33952 26140
rect 33976 26138 34032 26140
rect 33736 26086 33782 26138
rect 33782 26086 33792 26138
rect 33816 26086 33846 26138
rect 33846 26086 33858 26138
rect 33858 26086 33872 26138
rect 33896 26086 33910 26138
rect 33910 26086 33922 26138
rect 33922 26086 33952 26138
rect 33976 26086 33986 26138
rect 33986 26086 34032 26138
rect 33736 26084 33792 26086
rect 33816 26084 33872 26086
rect 33896 26084 33952 26086
rect 33976 26084 34032 26086
rect 2356 25594 2412 25596
rect 2436 25594 2492 25596
rect 2516 25594 2572 25596
rect 2596 25594 2652 25596
rect 2356 25542 2402 25594
rect 2402 25542 2412 25594
rect 2436 25542 2466 25594
rect 2466 25542 2478 25594
rect 2478 25542 2492 25594
rect 2516 25542 2530 25594
rect 2530 25542 2542 25594
rect 2542 25542 2572 25594
rect 2596 25542 2606 25594
rect 2606 25542 2652 25594
rect 2356 25540 2412 25542
rect 2436 25540 2492 25542
rect 2516 25540 2572 25542
rect 2596 25540 2652 25542
rect 33076 25594 33132 25596
rect 33156 25594 33212 25596
rect 33236 25594 33292 25596
rect 33316 25594 33372 25596
rect 33076 25542 33122 25594
rect 33122 25542 33132 25594
rect 33156 25542 33186 25594
rect 33186 25542 33198 25594
rect 33198 25542 33212 25594
rect 33236 25542 33250 25594
rect 33250 25542 33262 25594
rect 33262 25542 33292 25594
rect 33316 25542 33326 25594
rect 33326 25542 33372 25594
rect 33076 25540 33132 25542
rect 33156 25540 33212 25542
rect 33236 25540 33292 25542
rect 33316 25540 33372 25542
rect 3016 25050 3072 25052
rect 3096 25050 3152 25052
rect 3176 25050 3232 25052
rect 3256 25050 3312 25052
rect 3016 24998 3062 25050
rect 3062 24998 3072 25050
rect 3096 24998 3126 25050
rect 3126 24998 3138 25050
rect 3138 24998 3152 25050
rect 3176 24998 3190 25050
rect 3190 24998 3202 25050
rect 3202 24998 3232 25050
rect 3256 24998 3266 25050
rect 3266 24998 3312 25050
rect 3016 24996 3072 24998
rect 3096 24996 3152 24998
rect 3176 24996 3232 24998
rect 3256 24996 3312 24998
rect 33736 25050 33792 25052
rect 33816 25050 33872 25052
rect 33896 25050 33952 25052
rect 33976 25050 34032 25052
rect 33736 24998 33782 25050
rect 33782 24998 33792 25050
rect 33816 24998 33846 25050
rect 33846 24998 33858 25050
rect 33858 24998 33872 25050
rect 33896 24998 33910 25050
rect 33910 24998 33922 25050
rect 33922 24998 33952 25050
rect 33976 24998 33986 25050
rect 33986 24998 34032 25050
rect 33736 24996 33792 24998
rect 33816 24996 33872 24998
rect 33896 24996 33952 24998
rect 33976 24996 34032 24998
rect 2356 24506 2412 24508
rect 2436 24506 2492 24508
rect 2516 24506 2572 24508
rect 2596 24506 2652 24508
rect 2356 24454 2402 24506
rect 2402 24454 2412 24506
rect 2436 24454 2466 24506
rect 2466 24454 2478 24506
rect 2478 24454 2492 24506
rect 2516 24454 2530 24506
rect 2530 24454 2542 24506
rect 2542 24454 2572 24506
rect 2596 24454 2606 24506
rect 2606 24454 2652 24506
rect 2356 24452 2412 24454
rect 2436 24452 2492 24454
rect 2516 24452 2572 24454
rect 2596 24452 2652 24454
rect 33076 24506 33132 24508
rect 33156 24506 33212 24508
rect 33236 24506 33292 24508
rect 33316 24506 33372 24508
rect 33076 24454 33122 24506
rect 33122 24454 33132 24506
rect 33156 24454 33186 24506
rect 33186 24454 33198 24506
rect 33198 24454 33212 24506
rect 33236 24454 33250 24506
rect 33250 24454 33262 24506
rect 33262 24454 33292 24506
rect 33316 24454 33326 24506
rect 33326 24454 33372 24506
rect 33076 24452 33132 24454
rect 33156 24452 33212 24454
rect 33236 24452 33292 24454
rect 33316 24452 33372 24454
rect 3016 23962 3072 23964
rect 3096 23962 3152 23964
rect 3176 23962 3232 23964
rect 3256 23962 3312 23964
rect 3016 23910 3062 23962
rect 3062 23910 3072 23962
rect 3096 23910 3126 23962
rect 3126 23910 3138 23962
rect 3138 23910 3152 23962
rect 3176 23910 3190 23962
rect 3190 23910 3202 23962
rect 3202 23910 3232 23962
rect 3256 23910 3266 23962
rect 3266 23910 3312 23962
rect 3016 23908 3072 23910
rect 3096 23908 3152 23910
rect 3176 23908 3232 23910
rect 3256 23908 3312 23910
rect 33736 23962 33792 23964
rect 33816 23962 33872 23964
rect 33896 23962 33952 23964
rect 33976 23962 34032 23964
rect 33736 23910 33782 23962
rect 33782 23910 33792 23962
rect 33816 23910 33846 23962
rect 33846 23910 33858 23962
rect 33858 23910 33872 23962
rect 33896 23910 33910 23962
rect 33910 23910 33922 23962
rect 33922 23910 33952 23962
rect 33976 23910 33986 23962
rect 33986 23910 34032 23962
rect 33736 23908 33792 23910
rect 33816 23908 33872 23910
rect 33896 23908 33952 23910
rect 33976 23908 34032 23910
rect 2356 23418 2412 23420
rect 2436 23418 2492 23420
rect 2516 23418 2572 23420
rect 2596 23418 2652 23420
rect 2356 23366 2402 23418
rect 2402 23366 2412 23418
rect 2436 23366 2466 23418
rect 2466 23366 2478 23418
rect 2478 23366 2492 23418
rect 2516 23366 2530 23418
rect 2530 23366 2542 23418
rect 2542 23366 2572 23418
rect 2596 23366 2606 23418
rect 2606 23366 2652 23418
rect 2356 23364 2412 23366
rect 2436 23364 2492 23366
rect 2516 23364 2572 23366
rect 2596 23364 2652 23366
rect 33076 23418 33132 23420
rect 33156 23418 33212 23420
rect 33236 23418 33292 23420
rect 33316 23418 33372 23420
rect 33076 23366 33122 23418
rect 33122 23366 33132 23418
rect 33156 23366 33186 23418
rect 33186 23366 33198 23418
rect 33198 23366 33212 23418
rect 33236 23366 33250 23418
rect 33250 23366 33262 23418
rect 33262 23366 33292 23418
rect 33316 23366 33326 23418
rect 33326 23366 33372 23418
rect 33076 23364 33132 23366
rect 33156 23364 33212 23366
rect 33236 23364 33292 23366
rect 33316 23364 33372 23366
rect 3016 22874 3072 22876
rect 3096 22874 3152 22876
rect 3176 22874 3232 22876
rect 3256 22874 3312 22876
rect 3016 22822 3062 22874
rect 3062 22822 3072 22874
rect 3096 22822 3126 22874
rect 3126 22822 3138 22874
rect 3138 22822 3152 22874
rect 3176 22822 3190 22874
rect 3190 22822 3202 22874
rect 3202 22822 3232 22874
rect 3256 22822 3266 22874
rect 3266 22822 3312 22874
rect 3016 22820 3072 22822
rect 3096 22820 3152 22822
rect 3176 22820 3232 22822
rect 3256 22820 3312 22822
rect 33736 22874 33792 22876
rect 33816 22874 33872 22876
rect 33896 22874 33952 22876
rect 33976 22874 34032 22876
rect 33736 22822 33782 22874
rect 33782 22822 33792 22874
rect 33816 22822 33846 22874
rect 33846 22822 33858 22874
rect 33858 22822 33872 22874
rect 33896 22822 33910 22874
rect 33910 22822 33922 22874
rect 33922 22822 33952 22874
rect 33976 22822 33986 22874
rect 33986 22822 34032 22874
rect 33736 22820 33792 22822
rect 33816 22820 33872 22822
rect 33896 22820 33952 22822
rect 33976 22820 34032 22822
rect 2356 22330 2412 22332
rect 2436 22330 2492 22332
rect 2516 22330 2572 22332
rect 2596 22330 2652 22332
rect 2356 22278 2402 22330
rect 2402 22278 2412 22330
rect 2436 22278 2466 22330
rect 2466 22278 2478 22330
rect 2478 22278 2492 22330
rect 2516 22278 2530 22330
rect 2530 22278 2542 22330
rect 2542 22278 2572 22330
rect 2596 22278 2606 22330
rect 2606 22278 2652 22330
rect 2356 22276 2412 22278
rect 2436 22276 2492 22278
rect 2516 22276 2572 22278
rect 2596 22276 2652 22278
rect 33076 22330 33132 22332
rect 33156 22330 33212 22332
rect 33236 22330 33292 22332
rect 33316 22330 33372 22332
rect 33076 22278 33122 22330
rect 33122 22278 33132 22330
rect 33156 22278 33186 22330
rect 33186 22278 33198 22330
rect 33198 22278 33212 22330
rect 33236 22278 33250 22330
rect 33250 22278 33262 22330
rect 33262 22278 33292 22330
rect 33316 22278 33326 22330
rect 33326 22278 33372 22330
rect 33076 22276 33132 22278
rect 33156 22276 33212 22278
rect 33236 22276 33292 22278
rect 33316 22276 33372 22278
rect 3016 21786 3072 21788
rect 3096 21786 3152 21788
rect 3176 21786 3232 21788
rect 3256 21786 3312 21788
rect 3016 21734 3062 21786
rect 3062 21734 3072 21786
rect 3096 21734 3126 21786
rect 3126 21734 3138 21786
rect 3138 21734 3152 21786
rect 3176 21734 3190 21786
rect 3190 21734 3202 21786
rect 3202 21734 3232 21786
rect 3256 21734 3266 21786
rect 3266 21734 3312 21786
rect 3016 21732 3072 21734
rect 3096 21732 3152 21734
rect 3176 21732 3232 21734
rect 3256 21732 3312 21734
rect 33736 21786 33792 21788
rect 33816 21786 33872 21788
rect 33896 21786 33952 21788
rect 33976 21786 34032 21788
rect 33736 21734 33782 21786
rect 33782 21734 33792 21786
rect 33816 21734 33846 21786
rect 33846 21734 33858 21786
rect 33858 21734 33872 21786
rect 33896 21734 33910 21786
rect 33910 21734 33922 21786
rect 33922 21734 33952 21786
rect 33976 21734 33986 21786
rect 33986 21734 34032 21786
rect 33736 21732 33792 21734
rect 33816 21732 33872 21734
rect 33896 21732 33952 21734
rect 33976 21732 34032 21734
rect 2356 21242 2412 21244
rect 2436 21242 2492 21244
rect 2516 21242 2572 21244
rect 2596 21242 2652 21244
rect 2356 21190 2402 21242
rect 2402 21190 2412 21242
rect 2436 21190 2466 21242
rect 2466 21190 2478 21242
rect 2478 21190 2492 21242
rect 2516 21190 2530 21242
rect 2530 21190 2542 21242
rect 2542 21190 2572 21242
rect 2596 21190 2606 21242
rect 2606 21190 2652 21242
rect 2356 21188 2412 21190
rect 2436 21188 2492 21190
rect 2516 21188 2572 21190
rect 2596 21188 2652 21190
rect 33076 21242 33132 21244
rect 33156 21242 33212 21244
rect 33236 21242 33292 21244
rect 33316 21242 33372 21244
rect 33076 21190 33122 21242
rect 33122 21190 33132 21242
rect 33156 21190 33186 21242
rect 33186 21190 33198 21242
rect 33198 21190 33212 21242
rect 33236 21190 33250 21242
rect 33250 21190 33262 21242
rect 33262 21190 33292 21242
rect 33316 21190 33326 21242
rect 33326 21190 33372 21242
rect 33076 21188 33132 21190
rect 33156 21188 33212 21190
rect 33236 21188 33292 21190
rect 33316 21188 33372 21190
rect 3016 20698 3072 20700
rect 3096 20698 3152 20700
rect 3176 20698 3232 20700
rect 3256 20698 3312 20700
rect 3016 20646 3062 20698
rect 3062 20646 3072 20698
rect 3096 20646 3126 20698
rect 3126 20646 3138 20698
rect 3138 20646 3152 20698
rect 3176 20646 3190 20698
rect 3190 20646 3202 20698
rect 3202 20646 3232 20698
rect 3256 20646 3266 20698
rect 3266 20646 3312 20698
rect 3016 20644 3072 20646
rect 3096 20644 3152 20646
rect 3176 20644 3232 20646
rect 3256 20644 3312 20646
rect 33736 20698 33792 20700
rect 33816 20698 33872 20700
rect 33896 20698 33952 20700
rect 33976 20698 34032 20700
rect 33736 20646 33782 20698
rect 33782 20646 33792 20698
rect 33816 20646 33846 20698
rect 33846 20646 33858 20698
rect 33858 20646 33872 20698
rect 33896 20646 33910 20698
rect 33910 20646 33922 20698
rect 33922 20646 33952 20698
rect 33976 20646 33986 20698
rect 33986 20646 34032 20698
rect 33736 20644 33792 20646
rect 33816 20644 33872 20646
rect 33896 20644 33952 20646
rect 33976 20644 34032 20646
rect 2356 20154 2412 20156
rect 2436 20154 2492 20156
rect 2516 20154 2572 20156
rect 2596 20154 2652 20156
rect 2356 20102 2402 20154
rect 2402 20102 2412 20154
rect 2436 20102 2466 20154
rect 2466 20102 2478 20154
rect 2478 20102 2492 20154
rect 2516 20102 2530 20154
rect 2530 20102 2542 20154
rect 2542 20102 2572 20154
rect 2596 20102 2606 20154
rect 2606 20102 2652 20154
rect 2356 20100 2412 20102
rect 2436 20100 2492 20102
rect 2516 20100 2572 20102
rect 2596 20100 2652 20102
rect 33076 20154 33132 20156
rect 33156 20154 33212 20156
rect 33236 20154 33292 20156
rect 33316 20154 33372 20156
rect 33076 20102 33122 20154
rect 33122 20102 33132 20154
rect 33156 20102 33186 20154
rect 33186 20102 33198 20154
rect 33198 20102 33212 20154
rect 33236 20102 33250 20154
rect 33250 20102 33262 20154
rect 33262 20102 33292 20154
rect 33316 20102 33326 20154
rect 33326 20102 33372 20154
rect 33076 20100 33132 20102
rect 33156 20100 33212 20102
rect 33236 20100 33292 20102
rect 33316 20100 33372 20102
rect 3016 19610 3072 19612
rect 3096 19610 3152 19612
rect 3176 19610 3232 19612
rect 3256 19610 3312 19612
rect 3016 19558 3062 19610
rect 3062 19558 3072 19610
rect 3096 19558 3126 19610
rect 3126 19558 3138 19610
rect 3138 19558 3152 19610
rect 3176 19558 3190 19610
rect 3190 19558 3202 19610
rect 3202 19558 3232 19610
rect 3256 19558 3266 19610
rect 3266 19558 3312 19610
rect 3016 19556 3072 19558
rect 3096 19556 3152 19558
rect 3176 19556 3232 19558
rect 3256 19556 3312 19558
rect 33736 19610 33792 19612
rect 33816 19610 33872 19612
rect 33896 19610 33952 19612
rect 33976 19610 34032 19612
rect 33736 19558 33782 19610
rect 33782 19558 33792 19610
rect 33816 19558 33846 19610
rect 33846 19558 33858 19610
rect 33858 19558 33872 19610
rect 33896 19558 33910 19610
rect 33910 19558 33922 19610
rect 33922 19558 33952 19610
rect 33976 19558 33986 19610
rect 33986 19558 34032 19610
rect 33736 19556 33792 19558
rect 33816 19556 33872 19558
rect 33896 19556 33952 19558
rect 33976 19556 34032 19558
rect 2356 19066 2412 19068
rect 2436 19066 2492 19068
rect 2516 19066 2572 19068
rect 2596 19066 2652 19068
rect 2356 19014 2402 19066
rect 2402 19014 2412 19066
rect 2436 19014 2466 19066
rect 2466 19014 2478 19066
rect 2478 19014 2492 19066
rect 2516 19014 2530 19066
rect 2530 19014 2542 19066
rect 2542 19014 2572 19066
rect 2596 19014 2606 19066
rect 2606 19014 2652 19066
rect 2356 19012 2412 19014
rect 2436 19012 2492 19014
rect 2516 19012 2572 19014
rect 2596 19012 2652 19014
rect 33076 19066 33132 19068
rect 33156 19066 33212 19068
rect 33236 19066 33292 19068
rect 33316 19066 33372 19068
rect 33076 19014 33122 19066
rect 33122 19014 33132 19066
rect 33156 19014 33186 19066
rect 33186 19014 33198 19066
rect 33198 19014 33212 19066
rect 33236 19014 33250 19066
rect 33250 19014 33262 19066
rect 33262 19014 33292 19066
rect 33316 19014 33326 19066
rect 33326 19014 33372 19066
rect 33076 19012 33132 19014
rect 33156 19012 33212 19014
rect 33236 19012 33292 19014
rect 33316 19012 33372 19014
rect 3016 18522 3072 18524
rect 3096 18522 3152 18524
rect 3176 18522 3232 18524
rect 3256 18522 3312 18524
rect 3016 18470 3062 18522
rect 3062 18470 3072 18522
rect 3096 18470 3126 18522
rect 3126 18470 3138 18522
rect 3138 18470 3152 18522
rect 3176 18470 3190 18522
rect 3190 18470 3202 18522
rect 3202 18470 3232 18522
rect 3256 18470 3266 18522
rect 3266 18470 3312 18522
rect 3016 18468 3072 18470
rect 3096 18468 3152 18470
rect 3176 18468 3232 18470
rect 3256 18468 3312 18470
rect 33736 18522 33792 18524
rect 33816 18522 33872 18524
rect 33896 18522 33952 18524
rect 33976 18522 34032 18524
rect 33736 18470 33782 18522
rect 33782 18470 33792 18522
rect 33816 18470 33846 18522
rect 33846 18470 33858 18522
rect 33858 18470 33872 18522
rect 33896 18470 33910 18522
rect 33910 18470 33922 18522
rect 33922 18470 33952 18522
rect 33976 18470 33986 18522
rect 33986 18470 34032 18522
rect 33736 18468 33792 18470
rect 33816 18468 33872 18470
rect 33896 18468 33952 18470
rect 33976 18468 34032 18470
rect 2356 17978 2412 17980
rect 2436 17978 2492 17980
rect 2516 17978 2572 17980
rect 2596 17978 2652 17980
rect 2356 17926 2402 17978
rect 2402 17926 2412 17978
rect 2436 17926 2466 17978
rect 2466 17926 2478 17978
rect 2478 17926 2492 17978
rect 2516 17926 2530 17978
rect 2530 17926 2542 17978
rect 2542 17926 2572 17978
rect 2596 17926 2606 17978
rect 2606 17926 2652 17978
rect 2356 17924 2412 17926
rect 2436 17924 2492 17926
rect 2516 17924 2572 17926
rect 2596 17924 2652 17926
rect 33076 17978 33132 17980
rect 33156 17978 33212 17980
rect 33236 17978 33292 17980
rect 33316 17978 33372 17980
rect 33076 17926 33122 17978
rect 33122 17926 33132 17978
rect 33156 17926 33186 17978
rect 33186 17926 33198 17978
rect 33198 17926 33212 17978
rect 33236 17926 33250 17978
rect 33250 17926 33262 17978
rect 33262 17926 33292 17978
rect 33316 17926 33326 17978
rect 33326 17926 33372 17978
rect 33076 17924 33132 17926
rect 33156 17924 33212 17926
rect 33236 17924 33292 17926
rect 33316 17924 33372 17926
rect 3016 17434 3072 17436
rect 3096 17434 3152 17436
rect 3176 17434 3232 17436
rect 3256 17434 3312 17436
rect 3016 17382 3062 17434
rect 3062 17382 3072 17434
rect 3096 17382 3126 17434
rect 3126 17382 3138 17434
rect 3138 17382 3152 17434
rect 3176 17382 3190 17434
rect 3190 17382 3202 17434
rect 3202 17382 3232 17434
rect 3256 17382 3266 17434
rect 3266 17382 3312 17434
rect 3016 17380 3072 17382
rect 3096 17380 3152 17382
rect 3176 17380 3232 17382
rect 3256 17380 3312 17382
rect 33736 17434 33792 17436
rect 33816 17434 33872 17436
rect 33896 17434 33952 17436
rect 33976 17434 34032 17436
rect 33736 17382 33782 17434
rect 33782 17382 33792 17434
rect 33816 17382 33846 17434
rect 33846 17382 33858 17434
rect 33858 17382 33872 17434
rect 33896 17382 33910 17434
rect 33910 17382 33922 17434
rect 33922 17382 33952 17434
rect 33976 17382 33986 17434
rect 33986 17382 34032 17434
rect 33736 17380 33792 17382
rect 33816 17380 33872 17382
rect 33896 17380 33952 17382
rect 33976 17380 34032 17382
rect 2356 16890 2412 16892
rect 2436 16890 2492 16892
rect 2516 16890 2572 16892
rect 2596 16890 2652 16892
rect 2356 16838 2402 16890
rect 2402 16838 2412 16890
rect 2436 16838 2466 16890
rect 2466 16838 2478 16890
rect 2478 16838 2492 16890
rect 2516 16838 2530 16890
rect 2530 16838 2542 16890
rect 2542 16838 2572 16890
rect 2596 16838 2606 16890
rect 2606 16838 2652 16890
rect 2356 16836 2412 16838
rect 2436 16836 2492 16838
rect 2516 16836 2572 16838
rect 2596 16836 2652 16838
rect 33076 16890 33132 16892
rect 33156 16890 33212 16892
rect 33236 16890 33292 16892
rect 33316 16890 33372 16892
rect 33076 16838 33122 16890
rect 33122 16838 33132 16890
rect 33156 16838 33186 16890
rect 33186 16838 33198 16890
rect 33198 16838 33212 16890
rect 33236 16838 33250 16890
rect 33250 16838 33262 16890
rect 33262 16838 33292 16890
rect 33316 16838 33326 16890
rect 33326 16838 33372 16890
rect 33076 16836 33132 16838
rect 33156 16836 33212 16838
rect 33236 16836 33292 16838
rect 33316 16836 33372 16838
rect 3016 16346 3072 16348
rect 3096 16346 3152 16348
rect 3176 16346 3232 16348
rect 3256 16346 3312 16348
rect 3016 16294 3062 16346
rect 3062 16294 3072 16346
rect 3096 16294 3126 16346
rect 3126 16294 3138 16346
rect 3138 16294 3152 16346
rect 3176 16294 3190 16346
rect 3190 16294 3202 16346
rect 3202 16294 3232 16346
rect 3256 16294 3266 16346
rect 3266 16294 3312 16346
rect 3016 16292 3072 16294
rect 3096 16292 3152 16294
rect 3176 16292 3232 16294
rect 3256 16292 3312 16294
rect 33736 16346 33792 16348
rect 33816 16346 33872 16348
rect 33896 16346 33952 16348
rect 33976 16346 34032 16348
rect 33736 16294 33782 16346
rect 33782 16294 33792 16346
rect 33816 16294 33846 16346
rect 33846 16294 33858 16346
rect 33858 16294 33872 16346
rect 33896 16294 33910 16346
rect 33910 16294 33922 16346
rect 33922 16294 33952 16346
rect 33976 16294 33986 16346
rect 33986 16294 34032 16346
rect 33736 16292 33792 16294
rect 33816 16292 33872 16294
rect 33896 16292 33952 16294
rect 33976 16292 34032 16294
rect 2356 15802 2412 15804
rect 2436 15802 2492 15804
rect 2516 15802 2572 15804
rect 2596 15802 2652 15804
rect 2356 15750 2402 15802
rect 2402 15750 2412 15802
rect 2436 15750 2466 15802
rect 2466 15750 2478 15802
rect 2478 15750 2492 15802
rect 2516 15750 2530 15802
rect 2530 15750 2542 15802
rect 2542 15750 2572 15802
rect 2596 15750 2606 15802
rect 2606 15750 2652 15802
rect 2356 15748 2412 15750
rect 2436 15748 2492 15750
rect 2516 15748 2572 15750
rect 2596 15748 2652 15750
rect 33076 15802 33132 15804
rect 33156 15802 33212 15804
rect 33236 15802 33292 15804
rect 33316 15802 33372 15804
rect 33076 15750 33122 15802
rect 33122 15750 33132 15802
rect 33156 15750 33186 15802
rect 33186 15750 33198 15802
rect 33198 15750 33212 15802
rect 33236 15750 33250 15802
rect 33250 15750 33262 15802
rect 33262 15750 33292 15802
rect 33316 15750 33326 15802
rect 33326 15750 33372 15802
rect 33076 15748 33132 15750
rect 33156 15748 33212 15750
rect 33236 15748 33292 15750
rect 33316 15748 33372 15750
rect 3016 15258 3072 15260
rect 3096 15258 3152 15260
rect 3176 15258 3232 15260
rect 3256 15258 3312 15260
rect 3016 15206 3062 15258
rect 3062 15206 3072 15258
rect 3096 15206 3126 15258
rect 3126 15206 3138 15258
rect 3138 15206 3152 15258
rect 3176 15206 3190 15258
rect 3190 15206 3202 15258
rect 3202 15206 3232 15258
rect 3256 15206 3266 15258
rect 3266 15206 3312 15258
rect 3016 15204 3072 15206
rect 3096 15204 3152 15206
rect 3176 15204 3232 15206
rect 3256 15204 3312 15206
rect 33736 15258 33792 15260
rect 33816 15258 33872 15260
rect 33896 15258 33952 15260
rect 33976 15258 34032 15260
rect 33736 15206 33782 15258
rect 33782 15206 33792 15258
rect 33816 15206 33846 15258
rect 33846 15206 33858 15258
rect 33858 15206 33872 15258
rect 33896 15206 33910 15258
rect 33910 15206 33922 15258
rect 33922 15206 33952 15258
rect 33976 15206 33986 15258
rect 33986 15206 34032 15258
rect 33736 15204 33792 15206
rect 33816 15204 33872 15206
rect 33896 15204 33952 15206
rect 33976 15204 34032 15206
rect 58530 44920 58586 44976
rect 56506 15000 56562 15056
rect 2356 14714 2412 14716
rect 2436 14714 2492 14716
rect 2516 14714 2572 14716
rect 2596 14714 2652 14716
rect 2356 14662 2402 14714
rect 2402 14662 2412 14714
rect 2436 14662 2466 14714
rect 2466 14662 2478 14714
rect 2478 14662 2492 14714
rect 2516 14662 2530 14714
rect 2530 14662 2542 14714
rect 2542 14662 2572 14714
rect 2596 14662 2606 14714
rect 2606 14662 2652 14714
rect 2356 14660 2412 14662
rect 2436 14660 2492 14662
rect 2516 14660 2572 14662
rect 2596 14660 2652 14662
rect 33076 14714 33132 14716
rect 33156 14714 33212 14716
rect 33236 14714 33292 14716
rect 33316 14714 33372 14716
rect 33076 14662 33122 14714
rect 33122 14662 33132 14714
rect 33156 14662 33186 14714
rect 33186 14662 33198 14714
rect 33198 14662 33212 14714
rect 33236 14662 33250 14714
rect 33250 14662 33262 14714
rect 33262 14662 33292 14714
rect 33316 14662 33326 14714
rect 33326 14662 33372 14714
rect 33076 14660 33132 14662
rect 33156 14660 33212 14662
rect 33236 14660 33292 14662
rect 33316 14660 33372 14662
rect 3016 14170 3072 14172
rect 3096 14170 3152 14172
rect 3176 14170 3232 14172
rect 3256 14170 3312 14172
rect 3016 14118 3062 14170
rect 3062 14118 3072 14170
rect 3096 14118 3126 14170
rect 3126 14118 3138 14170
rect 3138 14118 3152 14170
rect 3176 14118 3190 14170
rect 3190 14118 3202 14170
rect 3202 14118 3232 14170
rect 3256 14118 3266 14170
rect 3266 14118 3312 14170
rect 3016 14116 3072 14118
rect 3096 14116 3152 14118
rect 3176 14116 3232 14118
rect 3256 14116 3312 14118
rect 33736 14170 33792 14172
rect 33816 14170 33872 14172
rect 33896 14170 33952 14172
rect 33976 14170 34032 14172
rect 33736 14118 33782 14170
rect 33782 14118 33792 14170
rect 33816 14118 33846 14170
rect 33846 14118 33858 14170
rect 33858 14118 33872 14170
rect 33896 14118 33910 14170
rect 33910 14118 33922 14170
rect 33922 14118 33952 14170
rect 33976 14118 33986 14170
rect 33986 14118 34032 14170
rect 33736 14116 33792 14118
rect 33816 14116 33872 14118
rect 33896 14116 33952 14118
rect 33976 14116 34032 14118
rect 2356 13626 2412 13628
rect 2436 13626 2492 13628
rect 2516 13626 2572 13628
rect 2596 13626 2652 13628
rect 2356 13574 2402 13626
rect 2402 13574 2412 13626
rect 2436 13574 2466 13626
rect 2466 13574 2478 13626
rect 2478 13574 2492 13626
rect 2516 13574 2530 13626
rect 2530 13574 2542 13626
rect 2542 13574 2572 13626
rect 2596 13574 2606 13626
rect 2606 13574 2652 13626
rect 2356 13572 2412 13574
rect 2436 13572 2492 13574
rect 2516 13572 2572 13574
rect 2596 13572 2652 13574
rect 33076 13626 33132 13628
rect 33156 13626 33212 13628
rect 33236 13626 33292 13628
rect 33316 13626 33372 13628
rect 33076 13574 33122 13626
rect 33122 13574 33132 13626
rect 33156 13574 33186 13626
rect 33186 13574 33198 13626
rect 33198 13574 33212 13626
rect 33236 13574 33250 13626
rect 33250 13574 33262 13626
rect 33262 13574 33292 13626
rect 33316 13574 33326 13626
rect 33326 13574 33372 13626
rect 33076 13572 33132 13574
rect 33156 13572 33212 13574
rect 33236 13572 33292 13574
rect 33316 13572 33372 13574
rect 3016 13082 3072 13084
rect 3096 13082 3152 13084
rect 3176 13082 3232 13084
rect 3256 13082 3312 13084
rect 3016 13030 3062 13082
rect 3062 13030 3072 13082
rect 3096 13030 3126 13082
rect 3126 13030 3138 13082
rect 3138 13030 3152 13082
rect 3176 13030 3190 13082
rect 3190 13030 3202 13082
rect 3202 13030 3232 13082
rect 3256 13030 3266 13082
rect 3266 13030 3312 13082
rect 3016 13028 3072 13030
rect 3096 13028 3152 13030
rect 3176 13028 3232 13030
rect 3256 13028 3312 13030
rect 33736 13082 33792 13084
rect 33816 13082 33872 13084
rect 33896 13082 33952 13084
rect 33976 13082 34032 13084
rect 33736 13030 33782 13082
rect 33782 13030 33792 13082
rect 33816 13030 33846 13082
rect 33846 13030 33858 13082
rect 33858 13030 33872 13082
rect 33896 13030 33910 13082
rect 33910 13030 33922 13082
rect 33922 13030 33952 13082
rect 33976 13030 33986 13082
rect 33986 13030 34032 13082
rect 33736 13028 33792 13030
rect 33816 13028 33872 13030
rect 33896 13028 33952 13030
rect 33976 13028 34032 13030
rect 2356 12538 2412 12540
rect 2436 12538 2492 12540
rect 2516 12538 2572 12540
rect 2596 12538 2652 12540
rect 2356 12486 2402 12538
rect 2402 12486 2412 12538
rect 2436 12486 2466 12538
rect 2466 12486 2478 12538
rect 2478 12486 2492 12538
rect 2516 12486 2530 12538
rect 2530 12486 2542 12538
rect 2542 12486 2572 12538
rect 2596 12486 2606 12538
rect 2606 12486 2652 12538
rect 2356 12484 2412 12486
rect 2436 12484 2492 12486
rect 2516 12484 2572 12486
rect 2596 12484 2652 12486
rect 33076 12538 33132 12540
rect 33156 12538 33212 12540
rect 33236 12538 33292 12540
rect 33316 12538 33372 12540
rect 33076 12486 33122 12538
rect 33122 12486 33132 12538
rect 33156 12486 33186 12538
rect 33186 12486 33198 12538
rect 33198 12486 33212 12538
rect 33236 12486 33250 12538
rect 33250 12486 33262 12538
rect 33262 12486 33292 12538
rect 33316 12486 33326 12538
rect 33326 12486 33372 12538
rect 33076 12484 33132 12486
rect 33156 12484 33212 12486
rect 33236 12484 33292 12486
rect 33316 12484 33372 12486
rect 3016 11994 3072 11996
rect 3096 11994 3152 11996
rect 3176 11994 3232 11996
rect 3256 11994 3312 11996
rect 3016 11942 3062 11994
rect 3062 11942 3072 11994
rect 3096 11942 3126 11994
rect 3126 11942 3138 11994
rect 3138 11942 3152 11994
rect 3176 11942 3190 11994
rect 3190 11942 3202 11994
rect 3202 11942 3232 11994
rect 3256 11942 3266 11994
rect 3266 11942 3312 11994
rect 3016 11940 3072 11942
rect 3096 11940 3152 11942
rect 3176 11940 3232 11942
rect 3256 11940 3312 11942
rect 33736 11994 33792 11996
rect 33816 11994 33872 11996
rect 33896 11994 33952 11996
rect 33976 11994 34032 11996
rect 33736 11942 33782 11994
rect 33782 11942 33792 11994
rect 33816 11942 33846 11994
rect 33846 11942 33858 11994
rect 33858 11942 33872 11994
rect 33896 11942 33910 11994
rect 33910 11942 33922 11994
rect 33922 11942 33952 11994
rect 33976 11942 33986 11994
rect 33986 11942 34032 11994
rect 33736 11940 33792 11942
rect 33816 11940 33872 11942
rect 33896 11940 33952 11942
rect 33976 11940 34032 11942
rect 2356 11450 2412 11452
rect 2436 11450 2492 11452
rect 2516 11450 2572 11452
rect 2596 11450 2652 11452
rect 2356 11398 2402 11450
rect 2402 11398 2412 11450
rect 2436 11398 2466 11450
rect 2466 11398 2478 11450
rect 2478 11398 2492 11450
rect 2516 11398 2530 11450
rect 2530 11398 2542 11450
rect 2542 11398 2572 11450
rect 2596 11398 2606 11450
rect 2606 11398 2652 11450
rect 2356 11396 2412 11398
rect 2436 11396 2492 11398
rect 2516 11396 2572 11398
rect 2596 11396 2652 11398
rect 33076 11450 33132 11452
rect 33156 11450 33212 11452
rect 33236 11450 33292 11452
rect 33316 11450 33372 11452
rect 33076 11398 33122 11450
rect 33122 11398 33132 11450
rect 33156 11398 33186 11450
rect 33186 11398 33198 11450
rect 33198 11398 33212 11450
rect 33236 11398 33250 11450
rect 33250 11398 33262 11450
rect 33262 11398 33292 11450
rect 33316 11398 33326 11450
rect 33326 11398 33372 11450
rect 33076 11396 33132 11398
rect 33156 11396 33212 11398
rect 33236 11396 33292 11398
rect 33316 11396 33372 11398
rect 3016 10906 3072 10908
rect 3096 10906 3152 10908
rect 3176 10906 3232 10908
rect 3256 10906 3312 10908
rect 3016 10854 3062 10906
rect 3062 10854 3072 10906
rect 3096 10854 3126 10906
rect 3126 10854 3138 10906
rect 3138 10854 3152 10906
rect 3176 10854 3190 10906
rect 3190 10854 3202 10906
rect 3202 10854 3232 10906
rect 3256 10854 3266 10906
rect 3266 10854 3312 10906
rect 3016 10852 3072 10854
rect 3096 10852 3152 10854
rect 3176 10852 3232 10854
rect 3256 10852 3312 10854
rect 33736 10906 33792 10908
rect 33816 10906 33872 10908
rect 33896 10906 33952 10908
rect 33976 10906 34032 10908
rect 33736 10854 33782 10906
rect 33782 10854 33792 10906
rect 33816 10854 33846 10906
rect 33846 10854 33858 10906
rect 33858 10854 33872 10906
rect 33896 10854 33910 10906
rect 33910 10854 33922 10906
rect 33922 10854 33952 10906
rect 33976 10854 33986 10906
rect 33986 10854 34032 10906
rect 33736 10852 33792 10854
rect 33816 10852 33872 10854
rect 33896 10852 33952 10854
rect 33976 10852 34032 10854
rect 2356 10362 2412 10364
rect 2436 10362 2492 10364
rect 2516 10362 2572 10364
rect 2596 10362 2652 10364
rect 2356 10310 2402 10362
rect 2402 10310 2412 10362
rect 2436 10310 2466 10362
rect 2466 10310 2478 10362
rect 2478 10310 2492 10362
rect 2516 10310 2530 10362
rect 2530 10310 2542 10362
rect 2542 10310 2572 10362
rect 2596 10310 2606 10362
rect 2606 10310 2652 10362
rect 2356 10308 2412 10310
rect 2436 10308 2492 10310
rect 2516 10308 2572 10310
rect 2596 10308 2652 10310
rect 33076 10362 33132 10364
rect 33156 10362 33212 10364
rect 33236 10362 33292 10364
rect 33316 10362 33372 10364
rect 33076 10310 33122 10362
rect 33122 10310 33132 10362
rect 33156 10310 33186 10362
rect 33186 10310 33198 10362
rect 33198 10310 33212 10362
rect 33236 10310 33250 10362
rect 33250 10310 33262 10362
rect 33262 10310 33292 10362
rect 33316 10310 33326 10362
rect 33326 10310 33372 10362
rect 33076 10308 33132 10310
rect 33156 10308 33212 10310
rect 33236 10308 33292 10310
rect 33316 10308 33372 10310
rect 3016 9818 3072 9820
rect 3096 9818 3152 9820
rect 3176 9818 3232 9820
rect 3256 9818 3312 9820
rect 3016 9766 3062 9818
rect 3062 9766 3072 9818
rect 3096 9766 3126 9818
rect 3126 9766 3138 9818
rect 3138 9766 3152 9818
rect 3176 9766 3190 9818
rect 3190 9766 3202 9818
rect 3202 9766 3232 9818
rect 3256 9766 3266 9818
rect 3266 9766 3312 9818
rect 3016 9764 3072 9766
rect 3096 9764 3152 9766
rect 3176 9764 3232 9766
rect 3256 9764 3312 9766
rect 33736 9818 33792 9820
rect 33816 9818 33872 9820
rect 33896 9818 33952 9820
rect 33976 9818 34032 9820
rect 33736 9766 33782 9818
rect 33782 9766 33792 9818
rect 33816 9766 33846 9818
rect 33846 9766 33858 9818
rect 33858 9766 33872 9818
rect 33896 9766 33910 9818
rect 33910 9766 33922 9818
rect 33922 9766 33952 9818
rect 33976 9766 33986 9818
rect 33986 9766 34032 9818
rect 33736 9764 33792 9766
rect 33816 9764 33872 9766
rect 33896 9764 33952 9766
rect 33976 9764 34032 9766
rect 2356 9274 2412 9276
rect 2436 9274 2492 9276
rect 2516 9274 2572 9276
rect 2596 9274 2652 9276
rect 2356 9222 2402 9274
rect 2402 9222 2412 9274
rect 2436 9222 2466 9274
rect 2466 9222 2478 9274
rect 2478 9222 2492 9274
rect 2516 9222 2530 9274
rect 2530 9222 2542 9274
rect 2542 9222 2572 9274
rect 2596 9222 2606 9274
rect 2606 9222 2652 9274
rect 2356 9220 2412 9222
rect 2436 9220 2492 9222
rect 2516 9220 2572 9222
rect 2596 9220 2652 9222
rect 33076 9274 33132 9276
rect 33156 9274 33212 9276
rect 33236 9274 33292 9276
rect 33316 9274 33372 9276
rect 33076 9222 33122 9274
rect 33122 9222 33132 9274
rect 33156 9222 33186 9274
rect 33186 9222 33198 9274
rect 33198 9222 33212 9274
rect 33236 9222 33250 9274
rect 33250 9222 33262 9274
rect 33262 9222 33292 9274
rect 33316 9222 33326 9274
rect 33326 9222 33372 9274
rect 33076 9220 33132 9222
rect 33156 9220 33212 9222
rect 33236 9220 33292 9222
rect 33316 9220 33372 9222
rect 3016 8730 3072 8732
rect 3096 8730 3152 8732
rect 3176 8730 3232 8732
rect 3256 8730 3312 8732
rect 3016 8678 3062 8730
rect 3062 8678 3072 8730
rect 3096 8678 3126 8730
rect 3126 8678 3138 8730
rect 3138 8678 3152 8730
rect 3176 8678 3190 8730
rect 3190 8678 3202 8730
rect 3202 8678 3232 8730
rect 3256 8678 3266 8730
rect 3266 8678 3312 8730
rect 3016 8676 3072 8678
rect 3096 8676 3152 8678
rect 3176 8676 3232 8678
rect 3256 8676 3312 8678
rect 33736 8730 33792 8732
rect 33816 8730 33872 8732
rect 33896 8730 33952 8732
rect 33976 8730 34032 8732
rect 33736 8678 33782 8730
rect 33782 8678 33792 8730
rect 33816 8678 33846 8730
rect 33846 8678 33858 8730
rect 33858 8678 33872 8730
rect 33896 8678 33910 8730
rect 33910 8678 33922 8730
rect 33922 8678 33952 8730
rect 33976 8678 33986 8730
rect 33986 8678 34032 8730
rect 33736 8676 33792 8678
rect 33816 8676 33872 8678
rect 33896 8676 33952 8678
rect 33976 8676 34032 8678
rect 2356 8186 2412 8188
rect 2436 8186 2492 8188
rect 2516 8186 2572 8188
rect 2596 8186 2652 8188
rect 2356 8134 2402 8186
rect 2402 8134 2412 8186
rect 2436 8134 2466 8186
rect 2466 8134 2478 8186
rect 2478 8134 2492 8186
rect 2516 8134 2530 8186
rect 2530 8134 2542 8186
rect 2542 8134 2572 8186
rect 2596 8134 2606 8186
rect 2606 8134 2652 8186
rect 2356 8132 2412 8134
rect 2436 8132 2492 8134
rect 2516 8132 2572 8134
rect 2596 8132 2652 8134
rect 33076 8186 33132 8188
rect 33156 8186 33212 8188
rect 33236 8186 33292 8188
rect 33316 8186 33372 8188
rect 33076 8134 33122 8186
rect 33122 8134 33132 8186
rect 33156 8134 33186 8186
rect 33186 8134 33198 8186
rect 33198 8134 33212 8186
rect 33236 8134 33250 8186
rect 33250 8134 33262 8186
rect 33262 8134 33292 8186
rect 33316 8134 33326 8186
rect 33326 8134 33372 8186
rect 33076 8132 33132 8134
rect 33156 8132 33212 8134
rect 33236 8132 33292 8134
rect 33316 8132 33372 8134
rect 3016 7642 3072 7644
rect 3096 7642 3152 7644
rect 3176 7642 3232 7644
rect 3256 7642 3312 7644
rect 3016 7590 3062 7642
rect 3062 7590 3072 7642
rect 3096 7590 3126 7642
rect 3126 7590 3138 7642
rect 3138 7590 3152 7642
rect 3176 7590 3190 7642
rect 3190 7590 3202 7642
rect 3202 7590 3232 7642
rect 3256 7590 3266 7642
rect 3266 7590 3312 7642
rect 3016 7588 3072 7590
rect 3096 7588 3152 7590
rect 3176 7588 3232 7590
rect 3256 7588 3312 7590
rect 33736 7642 33792 7644
rect 33816 7642 33872 7644
rect 33896 7642 33952 7644
rect 33976 7642 34032 7644
rect 33736 7590 33782 7642
rect 33782 7590 33792 7642
rect 33816 7590 33846 7642
rect 33846 7590 33858 7642
rect 33858 7590 33872 7642
rect 33896 7590 33910 7642
rect 33910 7590 33922 7642
rect 33922 7590 33952 7642
rect 33976 7590 33986 7642
rect 33986 7590 34032 7642
rect 33736 7588 33792 7590
rect 33816 7588 33872 7590
rect 33896 7588 33952 7590
rect 33976 7588 34032 7590
rect 2356 7098 2412 7100
rect 2436 7098 2492 7100
rect 2516 7098 2572 7100
rect 2596 7098 2652 7100
rect 2356 7046 2402 7098
rect 2402 7046 2412 7098
rect 2436 7046 2466 7098
rect 2466 7046 2478 7098
rect 2478 7046 2492 7098
rect 2516 7046 2530 7098
rect 2530 7046 2542 7098
rect 2542 7046 2572 7098
rect 2596 7046 2606 7098
rect 2606 7046 2652 7098
rect 2356 7044 2412 7046
rect 2436 7044 2492 7046
rect 2516 7044 2572 7046
rect 2596 7044 2652 7046
rect 33076 7098 33132 7100
rect 33156 7098 33212 7100
rect 33236 7098 33292 7100
rect 33316 7098 33372 7100
rect 33076 7046 33122 7098
rect 33122 7046 33132 7098
rect 33156 7046 33186 7098
rect 33186 7046 33198 7098
rect 33198 7046 33212 7098
rect 33236 7046 33250 7098
rect 33250 7046 33262 7098
rect 33262 7046 33292 7098
rect 33316 7046 33326 7098
rect 33326 7046 33372 7098
rect 33076 7044 33132 7046
rect 33156 7044 33212 7046
rect 33236 7044 33292 7046
rect 33316 7044 33372 7046
rect 3016 6554 3072 6556
rect 3096 6554 3152 6556
rect 3176 6554 3232 6556
rect 3256 6554 3312 6556
rect 3016 6502 3062 6554
rect 3062 6502 3072 6554
rect 3096 6502 3126 6554
rect 3126 6502 3138 6554
rect 3138 6502 3152 6554
rect 3176 6502 3190 6554
rect 3190 6502 3202 6554
rect 3202 6502 3232 6554
rect 3256 6502 3266 6554
rect 3266 6502 3312 6554
rect 3016 6500 3072 6502
rect 3096 6500 3152 6502
rect 3176 6500 3232 6502
rect 3256 6500 3312 6502
rect 33736 6554 33792 6556
rect 33816 6554 33872 6556
rect 33896 6554 33952 6556
rect 33976 6554 34032 6556
rect 33736 6502 33782 6554
rect 33782 6502 33792 6554
rect 33816 6502 33846 6554
rect 33846 6502 33858 6554
rect 33858 6502 33872 6554
rect 33896 6502 33910 6554
rect 33910 6502 33922 6554
rect 33922 6502 33952 6554
rect 33976 6502 33986 6554
rect 33986 6502 34032 6554
rect 33736 6500 33792 6502
rect 33816 6500 33872 6502
rect 33896 6500 33952 6502
rect 33976 6500 34032 6502
rect 2356 6010 2412 6012
rect 2436 6010 2492 6012
rect 2516 6010 2572 6012
rect 2596 6010 2652 6012
rect 2356 5958 2402 6010
rect 2402 5958 2412 6010
rect 2436 5958 2466 6010
rect 2466 5958 2478 6010
rect 2478 5958 2492 6010
rect 2516 5958 2530 6010
rect 2530 5958 2542 6010
rect 2542 5958 2572 6010
rect 2596 5958 2606 6010
rect 2606 5958 2652 6010
rect 2356 5956 2412 5958
rect 2436 5956 2492 5958
rect 2516 5956 2572 5958
rect 2596 5956 2652 5958
rect 33076 6010 33132 6012
rect 33156 6010 33212 6012
rect 33236 6010 33292 6012
rect 33316 6010 33372 6012
rect 33076 5958 33122 6010
rect 33122 5958 33132 6010
rect 33156 5958 33186 6010
rect 33186 5958 33198 6010
rect 33198 5958 33212 6010
rect 33236 5958 33250 6010
rect 33250 5958 33262 6010
rect 33262 5958 33292 6010
rect 33316 5958 33326 6010
rect 33326 5958 33372 6010
rect 33076 5956 33132 5958
rect 33156 5956 33212 5958
rect 33236 5956 33292 5958
rect 33316 5956 33372 5958
rect 3016 5466 3072 5468
rect 3096 5466 3152 5468
rect 3176 5466 3232 5468
rect 3256 5466 3312 5468
rect 3016 5414 3062 5466
rect 3062 5414 3072 5466
rect 3096 5414 3126 5466
rect 3126 5414 3138 5466
rect 3138 5414 3152 5466
rect 3176 5414 3190 5466
rect 3190 5414 3202 5466
rect 3202 5414 3232 5466
rect 3256 5414 3266 5466
rect 3266 5414 3312 5466
rect 3016 5412 3072 5414
rect 3096 5412 3152 5414
rect 3176 5412 3232 5414
rect 3256 5412 3312 5414
rect 33736 5466 33792 5468
rect 33816 5466 33872 5468
rect 33896 5466 33952 5468
rect 33976 5466 34032 5468
rect 33736 5414 33782 5466
rect 33782 5414 33792 5466
rect 33816 5414 33846 5466
rect 33846 5414 33858 5466
rect 33858 5414 33872 5466
rect 33896 5414 33910 5466
rect 33910 5414 33922 5466
rect 33922 5414 33952 5466
rect 33976 5414 33986 5466
rect 33986 5414 34032 5466
rect 33736 5412 33792 5414
rect 33816 5412 33872 5414
rect 33896 5412 33952 5414
rect 33976 5412 34032 5414
rect 2356 4922 2412 4924
rect 2436 4922 2492 4924
rect 2516 4922 2572 4924
rect 2596 4922 2652 4924
rect 2356 4870 2402 4922
rect 2402 4870 2412 4922
rect 2436 4870 2466 4922
rect 2466 4870 2478 4922
rect 2478 4870 2492 4922
rect 2516 4870 2530 4922
rect 2530 4870 2542 4922
rect 2542 4870 2572 4922
rect 2596 4870 2606 4922
rect 2606 4870 2652 4922
rect 2356 4868 2412 4870
rect 2436 4868 2492 4870
rect 2516 4868 2572 4870
rect 2596 4868 2652 4870
rect 33076 4922 33132 4924
rect 33156 4922 33212 4924
rect 33236 4922 33292 4924
rect 33316 4922 33372 4924
rect 33076 4870 33122 4922
rect 33122 4870 33132 4922
rect 33156 4870 33186 4922
rect 33186 4870 33198 4922
rect 33198 4870 33212 4922
rect 33236 4870 33250 4922
rect 33250 4870 33262 4922
rect 33262 4870 33292 4922
rect 33316 4870 33326 4922
rect 33326 4870 33372 4922
rect 33076 4868 33132 4870
rect 33156 4868 33212 4870
rect 33236 4868 33292 4870
rect 33316 4868 33372 4870
rect 3016 4378 3072 4380
rect 3096 4378 3152 4380
rect 3176 4378 3232 4380
rect 3256 4378 3312 4380
rect 3016 4326 3062 4378
rect 3062 4326 3072 4378
rect 3096 4326 3126 4378
rect 3126 4326 3138 4378
rect 3138 4326 3152 4378
rect 3176 4326 3190 4378
rect 3190 4326 3202 4378
rect 3202 4326 3232 4378
rect 3256 4326 3266 4378
rect 3266 4326 3312 4378
rect 3016 4324 3072 4326
rect 3096 4324 3152 4326
rect 3176 4324 3232 4326
rect 3256 4324 3312 4326
rect 33736 4378 33792 4380
rect 33816 4378 33872 4380
rect 33896 4378 33952 4380
rect 33976 4378 34032 4380
rect 33736 4326 33782 4378
rect 33782 4326 33792 4378
rect 33816 4326 33846 4378
rect 33846 4326 33858 4378
rect 33858 4326 33872 4378
rect 33896 4326 33910 4378
rect 33910 4326 33922 4378
rect 33922 4326 33952 4378
rect 33976 4326 33986 4378
rect 33986 4326 34032 4378
rect 33736 4324 33792 4326
rect 33816 4324 33872 4326
rect 33896 4324 33952 4326
rect 33976 4324 34032 4326
rect 2356 3834 2412 3836
rect 2436 3834 2492 3836
rect 2516 3834 2572 3836
rect 2596 3834 2652 3836
rect 2356 3782 2402 3834
rect 2402 3782 2412 3834
rect 2436 3782 2466 3834
rect 2466 3782 2478 3834
rect 2478 3782 2492 3834
rect 2516 3782 2530 3834
rect 2530 3782 2542 3834
rect 2542 3782 2572 3834
rect 2596 3782 2606 3834
rect 2606 3782 2652 3834
rect 2356 3780 2412 3782
rect 2436 3780 2492 3782
rect 2516 3780 2572 3782
rect 2596 3780 2652 3782
rect 33076 3834 33132 3836
rect 33156 3834 33212 3836
rect 33236 3834 33292 3836
rect 33316 3834 33372 3836
rect 33076 3782 33122 3834
rect 33122 3782 33132 3834
rect 33156 3782 33186 3834
rect 33186 3782 33198 3834
rect 33198 3782 33212 3834
rect 33236 3782 33250 3834
rect 33250 3782 33262 3834
rect 33262 3782 33292 3834
rect 33316 3782 33326 3834
rect 33326 3782 33372 3834
rect 33076 3780 33132 3782
rect 33156 3780 33212 3782
rect 33236 3780 33292 3782
rect 33316 3780 33372 3782
rect 3016 3290 3072 3292
rect 3096 3290 3152 3292
rect 3176 3290 3232 3292
rect 3256 3290 3312 3292
rect 3016 3238 3062 3290
rect 3062 3238 3072 3290
rect 3096 3238 3126 3290
rect 3126 3238 3138 3290
rect 3138 3238 3152 3290
rect 3176 3238 3190 3290
rect 3190 3238 3202 3290
rect 3202 3238 3232 3290
rect 3256 3238 3266 3290
rect 3266 3238 3312 3290
rect 3016 3236 3072 3238
rect 3096 3236 3152 3238
rect 3176 3236 3232 3238
rect 3256 3236 3312 3238
rect 33736 3290 33792 3292
rect 33816 3290 33872 3292
rect 33896 3290 33952 3292
rect 33976 3290 34032 3292
rect 33736 3238 33782 3290
rect 33782 3238 33792 3290
rect 33816 3238 33846 3290
rect 33846 3238 33858 3290
rect 33858 3238 33872 3290
rect 33896 3238 33910 3290
rect 33910 3238 33922 3290
rect 33922 3238 33952 3290
rect 33976 3238 33986 3290
rect 33986 3238 34032 3290
rect 33736 3236 33792 3238
rect 33816 3236 33872 3238
rect 33896 3236 33952 3238
rect 33976 3236 34032 3238
rect 2356 2746 2412 2748
rect 2436 2746 2492 2748
rect 2516 2746 2572 2748
rect 2596 2746 2652 2748
rect 2356 2694 2402 2746
rect 2402 2694 2412 2746
rect 2436 2694 2466 2746
rect 2466 2694 2478 2746
rect 2478 2694 2492 2746
rect 2516 2694 2530 2746
rect 2530 2694 2542 2746
rect 2542 2694 2572 2746
rect 2596 2694 2606 2746
rect 2606 2694 2652 2746
rect 2356 2692 2412 2694
rect 2436 2692 2492 2694
rect 2516 2692 2572 2694
rect 2596 2692 2652 2694
rect 33076 2746 33132 2748
rect 33156 2746 33212 2748
rect 33236 2746 33292 2748
rect 33316 2746 33372 2748
rect 33076 2694 33122 2746
rect 33122 2694 33132 2746
rect 33156 2694 33186 2746
rect 33186 2694 33198 2746
rect 33198 2694 33212 2746
rect 33236 2694 33250 2746
rect 33250 2694 33262 2746
rect 33262 2694 33292 2746
rect 33316 2694 33326 2746
rect 33326 2694 33372 2746
rect 33076 2692 33132 2694
rect 33156 2692 33212 2694
rect 33236 2692 33292 2694
rect 33316 2692 33372 2694
rect 3016 2202 3072 2204
rect 3096 2202 3152 2204
rect 3176 2202 3232 2204
rect 3256 2202 3312 2204
rect 3016 2150 3062 2202
rect 3062 2150 3072 2202
rect 3096 2150 3126 2202
rect 3126 2150 3138 2202
rect 3138 2150 3152 2202
rect 3176 2150 3190 2202
rect 3190 2150 3202 2202
rect 3202 2150 3232 2202
rect 3256 2150 3266 2202
rect 3266 2150 3312 2202
rect 3016 2148 3072 2150
rect 3096 2148 3152 2150
rect 3176 2148 3232 2150
rect 3256 2148 3312 2150
rect 33736 2202 33792 2204
rect 33816 2202 33872 2204
rect 33896 2202 33952 2204
rect 33976 2202 34032 2204
rect 33736 2150 33782 2202
rect 33782 2150 33792 2202
rect 33816 2150 33846 2202
rect 33846 2150 33858 2202
rect 33858 2150 33872 2202
rect 33896 2150 33910 2202
rect 33910 2150 33922 2202
rect 33922 2150 33952 2202
rect 33976 2150 33986 2202
rect 33986 2150 34032 2202
rect 33736 2148 33792 2150
rect 33816 2148 33872 2150
rect 33896 2148 33952 2150
rect 33976 2148 34032 2150
<< metal3 >>
rect 3006 57696 3322 57697
rect 3006 57632 3012 57696
rect 3076 57632 3092 57696
rect 3156 57632 3172 57696
rect 3236 57632 3252 57696
rect 3316 57632 3322 57696
rect 3006 57631 3322 57632
rect 33726 57696 34042 57697
rect 33726 57632 33732 57696
rect 33796 57632 33812 57696
rect 33876 57632 33892 57696
rect 33956 57632 33972 57696
rect 34036 57632 34042 57696
rect 33726 57631 34042 57632
rect 2346 57152 2662 57153
rect 2346 57088 2352 57152
rect 2416 57088 2432 57152
rect 2496 57088 2512 57152
rect 2576 57088 2592 57152
rect 2656 57088 2662 57152
rect 2346 57087 2662 57088
rect 33066 57152 33382 57153
rect 33066 57088 33072 57152
rect 33136 57088 33152 57152
rect 33216 57088 33232 57152
rect 33296 57088 33312 57152
rect 33376 57088 33382 57152
rect 33066 57087 33382 57088
rect 3006 56608 3322 56609
rect 3006 56544 3012 56608
rect 3076 56544 3092 56608
rect 3156 56544 3172 56608
rect 3236 56544 3252 56608
rect 3316 56544 3322 56608
rect 3006 56543 3322 56544
rect 33726 56608 34042 56609
rect 33726 56544 33732 56608
rect 33796 56544 33812 56608
rect 33876 56544 33892 56608
rect 33956 56544 33972 56608
rect 34036 56544 34042 56608
rect 33726 56543 34042 56544
rect 17401 56538 17467 56541
rect 19885 56538 19951 56541
rect 17401 56536 19951 56538
rect 17401 56480 17406 56536
rect 17462 56480 19890 56536
rect 19946 56480 19951 56536
rect 17401 56478 19951 56480
rect 17401 56475 17467 56478
rect 19885 56475 19951 56478
rect 2346 56064 2662 56065
rect 2346 56000 2352 56064
rect 2416 56000 2432 56064
rect 2496 56000 2512 56064
rect 2576 56000 2592 56064
rect 2656 56000 2662 56064
rect 2346 55999 2662 56000
rect 33066 56064 33382 56065
rect 33066 56000 33072 56064
rect 33136 56000 33152 56064
rect 33216 56000 33232 56064
rect 33296 56000 33312 56064
rect 33376 56000 33382 56064
rect 33066 55999 33382 56000
rect 20529 55858 20595 55861
rect 21909 55858 21975 55861
rect 20529 55856 21975 55858
rect 20529 55800 20534 55856
rect 20590 55800 21914 55856
rect 21970 55800 21975 55856
rect 20529 55798 21975 55800
rect 20529 55795 20595 55798
rect 21909 55795 21975 55798
rect 17217 55586 17283 55589
rect 19609 55586 19675 55589
rect 22829 55586 22895 55589
rect 17217 55584 22895 55586
rect 17217 55528 17222 55584
rect 17278 55528 19614 55584
rect 19670 55528 22834 55584
rect 22890 55528 22895 55584
rect 17217 55526 22895 55528
rect 17217 55523 17283 55526
rect 19609 55523 19675 55526
rect 22829 55523 22895 55526
rect 3006 55520 3322 55521
rect 3006 55456 3012 55520
rect 3076 55456 3092 55520
rect 3156 55456 3172 55520
rect 3236 55456 3252 55520
rect 3316 55456 3322 55520
rect 3006 55455 3322 55456
rect 33726 55520 34042 55521
rect 33726 55456 33732 55520
rect 33796 55456 33812 55520
rect 33876 55456 33892 55520
rect 33956 55456 33972 55520
rect 34036 55456 34042 55520
rect 33726 55455 34042 55456
rect 16941 55314 17007 55317
rect 17309 55314 17375 55317
rect 49049 55314 49115 55317
rect 16941 55312 49115 55314
rect 16941 55256 16946 55312
rect 17002 55256 17314 55312
rect 17370 55256 49054 55312
rect 49110 55256 49115 55312
rect 16941 55254 49115 55256
rect 16941 55251 17007 55254
rect 17309 55251 17375 55254
rect 49049 55251 49115 55254
rect 2346 54976 2662 54977
rect 2346 54912 2352 54976
rect 2416 54912 2432 54976
rect 2496 54912 2512 54976
rect 2576 54912 2592 54976
rect 2656 54912 2662 54976
rect 2346 54911 2662 54912
rect 33066 54976 33382 54977
rect 33066 54912 33072 54976
rect 33136 54912 33152 54976
rect 33216 54912 33232 54976
rect 33296 54912 33312 54976
rect 33376 54912 33382 54976
rect 33066 54911 33382 54912
rect 3006 54432 3322 54433
rect 3006 54368 3012 54432
rect 3076 54368 3092 54432
rect 3156 54368 3172 54432
rect 3236 54368 3252 54432
rect 3316 54368 3322 54432
rect 3006 54367 3322 54368
rect 33726 54432 34042 54433
rect 33726 54368 33732 54432
rect 33796 54368 33812 54432
rect 33876 54368 33892 54432
rect 33956 54368 33972 54432
rect 34036 54368 34042 54432
rect 33726 54367 34042 54368
rect 2346 53888 2662 53889
rect 2346 53824 2352 53888
rect 2416 53824 2432 53888
rect 2496 53824 2512 53888
rect 2576 53824 2592 53888
rect 2656 53824 2662 53888
rect 2346 53823 2662 53824
rect 33066 53888 33382 53889
rect 33066 53824 33072 53888
rect 33136 53824 33152 53888
rect 33216 53824 33232 53888
rect 33296 53824 33312 53888
rect 33376 53824 33382 53888
rect 33066 53823 33382 53824
rect 3006 53344 3322 53345
rect 3006 53280 3012 53344
rect 3076 53280 3092 53344
rect 3156 53280 3172 53344
rect 3236 53280 3252 53344
rect 3316 53280 3322 53344
rect 3006 53279 3322 53280
rect 33726 53344 34042 53345
rect 33726 53280 33732 53344
rect 33796 53280 33812 53344
rect 33876 53280 33892 53344
rect 33956 53280 33972 53344
rect 34036 53280 34042 53344
rect 33726 53279 34042 53280
rect 2346 52800 2662 52801
rect 2346 52736 2352 52800
rect 2416 52736 2432 52800
rect 2496 52736 2512 52800
rect 2576 52736 2592 52800
rect 2656 52736 2662 52800
rect 2346 52735 2662 52736
rect 33066 52800 33382 52801
rect 33066 52736 33072 52800
rect 33136 52736 33152 52800
rect 33216 52736 33232 52800
rect 33296 52736 33312 52800
rect 33376 52736 33382 52800
rect 33066 52735 33382 52736
rect 3006 52256 3322 52257
rect 3006 52192 3012 52256
rect 3076 52192 3092 52256
rect 3156 52192 3172 52256
rect 3236 52192 3252 52256
rect 3316 52192 3322 52256
rect 3006 52191 3322 52192
rect 33726 52256 34042 52257
rect 33726 52192 33732 52256
rect 33796 52192 33812 52256
rect 33876 52192 33892 52256
rect 33956 52192 33972 52256
rect 34036 52192 34042 52256
rect 33726 52191 34042 52192
rect 2346 51712 2662 51713
rect 2346 51648 2352 51712
rect 2416 51648 2432 51712
rect 2496 51648 2512 51712
rect 2576 51648 2592 51712
rect 2656 51648 2662 51712
rect 2346 51647 2662 51648
rect 33066 51712 33382 51713
rect 33066 51648 33072 51712
rect 33136 51648 33152 51712
rect 33216 51648 33232 51712
rect 33296 51648 33312 51712
rect 33376 51648 33382 51712
rect 33066 51647 33382 51648
rect 3006 51168 3322 51169
rect 3006 51104 3012 51168
rect 3076 51104 3092 51168
rect 3156 51104 3172 51168
rect 3236 51104 3252 51168
rect 3316 51104 3322 51168
rect 3006 51103 3322 51104
rect 33726 51168 34042 51169
rect 33726 51104 33732 51168
rect 33796 51104 33812 51168
rect 33876 51104 33892 51168
rect 33956 51104 33972 51168
rect 34036 51104 34042 51168
rect 33726 51103 34042 51104
rect 2346 50624 2662 50625
rect 2346 50560 2352 50624
rect 2416 50560 2432 50624
rect 2496 50560 2512 50624
rect 2576 50560 2592 50624
rect 2656 50560 2662 50624
rect 2346 50559 2662 50560
rect 33066 50624 33382 50625
rect 33066 50560 33072 50624
rect 33136 50560 33152 50624
rect 33216 50560 33232 50624
rect 33296 50560 33312 50624
rect 33376 50560 33382 50624
rect 33066 50559 33382 50560
rect 3006 50080 3322 50081
rect 3006 50016 3012 50080
rect 3076 50016 3092 50080
rect 3156 50016 3172 50080
rect 3236 50016 3252 50080
rect 3316 50016 3322 50080
rect 3006 50015 3322 50016
rect 33726 50080 34042 50081
rect 33726 50016 33732 50080
rect 33796 50016 33812 50080
rect 33876 50016 33892 50080
rect 33956 50016 33972 50080
rect 34036 50016 34042 50080
rect 33726 50015 34042 50016
rect 2346 49536 2662 49537
rect 2346 49472 2352 49536
rect 2416 49472 2432 49536
rect 2496 49472 2512 49536
rect 2576 49472 2592 49536
rect 2656 49472 2662 49536
rect 2346 49471 2662 49472
rect 33066 49536 33382 49537
rect 33066 49472 33072 49536
rect 33136 49472 33152 49536
rect 33216 49472 33232 49536
rect 33296 49472 33312 49536
rect 33376 49472 33382 49536
rect 33066 49471 33382 49472
rect 3006 48992 3322 48993
rect 3006 48928 3012 48992
rect 3076 48928 3092 48992
rect 3156 48928 3172 48992
rect 3236 48928 3252 48992
rect 3316 48928 3322 48992
rect 3006 48927 3322 48928
rect 33726 48992 34042 48993
rect 33726 48928 33732 48992
rect 33796 48928 33812 48992
rect 33876 48928 33892 48992
rect 33956 48928 33972 48992
rect 34036 48928 34042 48992
rect 33726 48927 34042 48928
rect 2346 48448 2662 48449
rect 2346 48384 2352 48448
rect 2416 48384 2432 48448
rect 2496 48384 2512 48448
rect 2576 48384 2592 48448
rect 2656 48384 2662 48448
rect 2346 48383 2662 48384
rect 33066 48448 33382 48449
rect 33066 48384 33072 48448
rect 33136 48384 33152 48448
rect 33216 48384 33232 48448
rect 33296 48384 33312 48448
rect 33376 48384 33382 48448
rect 33066 48383 33382 48384
rect 3006 47904 3322 47905
rect 3006 47840 3012 47904
rect 3076 47840 3092 47904
rect 3156 47840 3172 47904
rect 3236 47840 3252 47904
rect 3316 47840 3322 47904
rect 3006 47839 3322 47840
rect 33726 47904 34042 47905
rect 33726 47840 33732 47904
rect 33796 47840 33812 47904
rect 33876 47840 33892 47904
rect 33956 47840 33972 47904
rect 34036 47840 34042 47904
rect 33726 47839 34042 47840
rect 2346 47360 2662 47361
rect 2346 47296 2352 47360
rect 2416 47296 2432 47360
rect 2496 47296 2512 47360
rect 2576 47296 2592 47360
rect 2656 47296 2662 47360
rect 2346 47295 2662 47296
rect 33066 47360 33382 47361
rect 33066 47296 33072 47360
rect 33136 47296 33152 47360
rect 33216 47296 33232 47360
rect 33296 47296 33312 47360
rect 33376 47296 33382 47360
rect 33066 47295 33382 47296
rect 3006 46816 3322 46817
rect 3006 46752 3012 46816
rect 3076 46752 3092 46816
rect 3156 46752 3172 46816
rect 3236 46752 3252 46816
rect 3316 46752 3322 46816
rect 3006 46751 3322 46752
rect 33726 46816 34042 46817
rect 33726 46752 33732 46816
rect 33796 46752 33812 46816
rect 33876 46752 33892 46816
rect 33956 46752 33972 46816
rect 34036 46752 34042 46816
rect 33726 46751 34042 46752
rect 2346 46272 2662 46273
rect 2346 46208 2352 46272
rect 2416 46208 2432 46272
rect 2496 46208 2512 46272
rect 2576 46208 2592 46272
rect 2656 46208 2662 46272
rect 2346 46207 2662 46208
rect 33066 46272 33382 46273
rect 33066 46208 33072 46272
rect 33136 46208 33152 46272
rect 33216 46208 33232 46272
rect 33296 46208 33312 46272
rect 33376 46208 33382 46272
rect 33066 46207 33382 46208
rect 3006 45728 3322 45729
rect 3006 45664 3012 45728
rect 3076 45664 3092 45728
rect 3156 45664 3172 45728
rect 3236 45664 3252 45728
rect 3316 45664 3322 45728
rect 3006 45663 3322 45664
rect 33726 45728 34042 45729
rect 33726 45664 33732 45728
rect 33796 45664 33812 45728
rect 33876 45664 33892 45728
rect 33956 45664 33972 45728
rect 34036 45664 34042 45728
rect 33726 45663 34042 45664
rect 2346 45184 2662 45185
rect 2346 45120 2352 45184
rect 2416 45120 2432 45184
rect 2496 45120 2512 45184
rect 2576 45120 2592 45184
rect 2656 45120 2662 45184
rect 2346 45119 2662 45120
rect 33066 45184 33382 45185
rect 33066 45120 33072 45184
rect 33136 45120 33152 45184
rect 33216 45120 33232 45184
rect 33296 45120 33312 45184
rect 33376 45120 33382 45184
rect 33066 45119 33382 45120
rect 58525 44978 58591 44981
rect 59200 44978 60000 45008
rect 58525 44976 60000 44978
rect 58525 44920 58530 44976
rect 58586 44920 60000 44976
rect 58525 44918 60000 44920
rect 58525 44915 58591 44918
rect 59200 44888 60000 44918
rect 3006 44640 3322 44641
rect 3006 44576 3012 44640
rect 3076 44576 3092 44640
rect 3156 44576 3172 44640
rect 3236 44576 3252 44640
rect 3316 44576 3322 44640
rect 3006 44575 3322 44576
rect 33726 44640 34042 44641
rect 33726 44576 33732 44640
rect 33796 44576 33812 44640
rect 33876 44576 33892 44640
rect 33956 44576 33972 44640
rect 34036 44576 34042 44640
rect 33726 44575 34042 44576
rect 2346 44096 2662 44097
rect 2346 44032 2352 44096
rect 2416 44032 2432 44096
rect 2496 44032 2512 44096
rect 2576 44032 2592 44096
rect 2656 44032 2662 44096
rect 2346 44031 2662 44032
rect 33066 44096 33382 44097
rect 33066 44032 33072 44096
rect 33136 44032 33152 44096
rect 33216 44032 33232 44096
rect 33296 44032 33312 44096
rect 33376 44032 33382 44096
rect 33066 44031 33382 44032
rect 3006 43552 3322 43553
rect 3006 43488 3012 43552
rect 3076 43488 3092 43552
rect 3156 43488 3172 43552
rect 3236 43488 3252 43552
rect 3316 43488 3322 43552
rect 3006 43487 3322 43488
rect 33726 43552 34042 43553
rect 33726 43488 33732 43552
rect 33796 43488 33812 43552
rect 33876 43488 33892 43552
rect 33956 43488 33972 43552
rect 34036 43488 34042 43552
rect 33726 43487 34042 43488
rect 2346 43008 2662 43009
rect 2346 42944 2352 43008
rect 2416 42944 2432 43008
rect 2496 42944 2512 43008
rect 2576 42944 2592 43008
rect 2656 42944 2662 43008
rect 2346 42943 2662 42944
rect 33066 43008 33382 43009
rect 33066 42944 33072 43008
rect 33136 42944 33152 43008
rect 33216 42944 33232 43008
rect 33296 42944 33312 43008
rect 33376 42944 33382 43008
rect 33066 42943 33382 42944
rect 3006 42464 3322 42465
rect 3006 42400 3012 42464
rect 3076 42400 3092 42464
rect 3156 42400 3172 42464
rect 3236 42400 3252 42464
rect 3316 42400 3322 42464
rect 3006 42399 3322 42400
rect 33726 42464 34042 42465
rect 33726 42400 33732 42464
rect 33796 42400 33812 42464
rect 33876 42400 33892 42464
rect 33956 42400 33972 42464
rect 34036 42400 34042 42464
rect 33726 42399 34042 42400
rect 2346 41920 2662 41921
rect 2346 41856 2352 41920
rect 2416 41856 2432 41920
rect 2496 41856 2512 41920
rect 2576 41856 2592 41920
rect 2656 41856 2662 41920
rect 2346 41855 2662 41856
rect 33066 41920 33382 41921
rect 33066 41856 33072 41920
rect 33136 41856 33152 41920
rect 33216 41856 33232 41920
rect 33296 41856 33312 41920
rect 33376 41856 33382 41920
rect 33066 41855 33382 41856
rect 3006 41376 3322 41377
rect 3006 41312 3012 41376
rect 3076 41312 3092 41376
rect 3156 41312 3172 41376
rect 3236 41312 3252 41376
rect 3316 41312 3322 41376
rect 3006 41311 3322 41312
rect 33726 41376 34042 41377
rect 33726 41312 33732 41376
rect 33796 41312 33812 41376
rect 33876 41312 33892 41376
rect 33956 41312 33972 41376
rect 34036 41312 34042 41376
rect 33726 41311 34042 41312
rect 2346 40832 2662 40833
rect 2346 40768 2352 40832
rect 2416 40768 2432 40832
rect 2496 40768 2512 40832
rect 2576 40768 2592 40832
rect 2656 40768 2662 40832
rect 2346 40767 2662 40768
rect 33066 40832 33382 40833
rect 33066 40768 33072 40832
rect 33136 40768 33152 40832
rect 33216 40768 33232 40832
rect 33296 40768 33312 40832
rect 33376 40768 33382 40832
rect 33066 40767 33382 40768
rect 3006 40288 3322 40289
rect 3006 40224 3012 40288
rect 3076 40224 3092 40288
rect 3156 40224 3172 40288
rect 3236 40224 3252 40288
rect 3316 40224 3322 40288
rect 3006 40223 3322 40224
rect 33726 40288 34042 40289
rect 33726 40224 33732 40288
rect 33796 40224 33812 40288
rect 33876 40224 33892 40288
rect 33956 40224 33972 40288
rect 34036 40224 34042 40288
rect 33726 40223 34042 40224
rect 2346 39744 2662 39745
rect 2346 39680 2352 39744
rect 2416 39680 2432 39744
rect 2496 39680 2512 39744
rect 2576 39680 2592 39744
rect 2656 39680 2662 39744
rect 2346 39679 2662 39680
rect 33066 39744 33382 39745
rect 33066 39680 33072 39744
rect 33136 39680 33152 39744
rect 33216 39680 33232 39744
rect 33296 39680 33312 39744
rect 33376 39680 33382 39744
rect 33066 39679 33382 39680
rect 3006 39200 3322 39201
rect 3006 39136 3012 39200
rect 3076 39136 3092 39200
rect 3156 39136 3172 39200
rect 3236 39136 3252 39200
rect 3316 39136 3322 39200
rect 3006 39135 3322 39136
rect 33726 39200 34042 39201
rect 33726 39136 33732 39200
rect 33796 39136 33812 39200
rect 33876 39136 33892 39200
rect 33956 39136 33972 39200
rect 34036 39136 34042 39200
rect 33726 39135 34042 39136
rect 2346 38656 2662 38657
rect 2346 38592 2352 38656
rect 2416 38592 2432 38656
rect 2496 38592 2512 38656
rect 2576 38592 2592 38656
rect 2656 38592 2662 38656
rect 2346 38591 2662 38592
rect 33066 38656 33382 38657
rect 33066 38592 33072 38656
rect 33136 38592 33152 38656
rect 33216 38592 33232 38656
rect 33296 38592 33312 38656
rect 33376 38592 33382 38656
rect 33066 38591 33382 38592
rect 3006 38112 3322 38113
rect 3006 38048 3012 38112
rect 3076 38048 3092 38112
rect 3156 38048 3172 38112
rect 3236 38048 3252 38112
rect 3316 38048 3322 38112
rect 3006 38047 3322 38048
rect 33726 38112 34042 38113
rect 33726 38048 33732 38112
rect 33796 38048 33812 38112
rect 33876 38048 33892 38112
rect 33956 38048 33972 38112
rect 34036 38048 34042 38112
rect 33726 38047 34042 38048
rect 2346 37568 2662 37569
rect 2346 37504 2352 37568
rect 2416 37504 2432 37568
rect 2496 37504 2512 37568
rect 2576 37504 2592 37568
rect 2656 37504 2662 37568
rect 2346 37503 2662 37504
rect 33066 37568 33382 37569
rect 33066 37504 33072 37568
rect 33136 37504 33152 37568
rect 33216 37504 33232 37568
rect 33296 37504 33312 37568
rect 33376 37504 33382 37568
rect 33066 37503 33382 37504
rect 3006 37024 3322 37025
rect 3006 36960 3012 37024
rect 3076 36960 3092 37024
rect 3156 36960 3172 37024
rect 3236 36960 3252 37024
rect 3316 36960 3322 37024
rect 3006 36959 3322 36960
rect 33726 37024 34042 37025
rect 33726 36960 33732 37024
rect 33796 36960 33812 37024
rect 33876 36960 33892 37024
rect 33956 36960 33972 37024
rect 34036 36960 34042 37024
rect 33726 36959 34042 36960
rect 2346 36480 2662 36481
rect 2346 36416 2352 36480
rect 2416 36416 2432 36480
rect 2496 36416 2512 36480
rect 2576 36416 2592 36480
rect 2656 36416 2662 36480
rect 2346 36415 2662 36416
rect 33066 36480 33382 36481
rect 33066 36416 33072 36480
rect 33136 36416 33152 36480
rect 33216 36416 33232 36480
rect 33296 36416 33312 36480
rect 33376 36416 33382 36480
rect 33066 36415 33382 36416
rect 3006 35936 3322 35937
rect 3006 35872 3012 35936
rect 3076 35872 3092 35936
rect 3156 35872 3172 35936
rect 3236 35872 3252 35936
rect 3316 35872 3322 35936
rect 3006 35871 3322 35872
rect 33726 35936 34042 35937
rect 33726 35872 33732 35936
rect 33796 35872 33812 35936
rect 33876 35872 33892 35936
rect 33956 35872 33972 35936
rect 34036 35872 34042 35936
rect 33726 35871 34042 35872
rect 2346 35392 2662 35393
rect 2346 35328 2352 35392
rect 2416 35328 2432 35392
rect 2496 35328 2512 35392
rect 2576 35328 2592 35392
rect 2656 35328 2662 35392
rect 2346 35327 2662 35328
rect 33066 35392 33382 35393
rect 33066 35328 33072 35392
rect 33136 35328 33152 35392
rect 33216 35328 33232 35392
rect 33296 35328 33312 35392
rect 33376 35328 33382 35392
rect 33066 35327 33382 35328
rect 3006 34848 3322 34849
rect 3006 34784 3012 34848
rect 3076 34784 3092 34848
rect 3156 34784 3172 34848
rect 3236 34784 3252 34848
rect 3316 34784 3322 34848
rect 3006 34783 3322 34784
rect 33726 34848 34042 34849
rect 33726 34784 33732 34848
rect 33796 34784 33812 34848
rect 33876 34784 33892 34848
rect 33956 34784 33972 34848
rect 34036 34784 34042 34848
rect 33726 34783 34042 34784
rect 2346 34304 2662 34305
rect 2346 34240 2352 34304
rect 2416 34240 2432 34304
rect 2496 34240 2512 34304
rect 2576 34240 2592 34304
rect 2656 34240 2662 34304
rect 2346 34239 2662 34240
rect 33066 34304 33382 34305
rect 33066 34240 33072 34304
rect 33136 34240 33152 34304
rect 33216 34240 33232 34304
rect 33296 34240 33312 34304
rect 33376 34240 33382 34304
rect 33066 34239 33382 34240
rect 3006 33760 3322 33761
rect 3006 33696 3012 33760
rect 3076 33696 3092 33760
rect 3156 33696 3172 33760
rect 3236 33696 3252 33760
rect 3316 33696 3322 33760
rect 3006 33695 3322 33696
rect 33726 33760 34042 33761
rect 33726 33696 33732 33760
rect 33796 33696 33812 33760
rect 33876 33696 33892 33760
rect 33956 33696 33972 33760
rect 34036 33696 34042 33760
rect 33726 33695 34042 33696
rect 2346 33216 2662 33217
rect 2346 33152 2352 33216
rect 2416 33152 2432 33216
rect 2496 33152 2512 33216
rect 2576 33152 2592 33216
rect 2656 33152 2662 33216
rect 2346 33151 2662 33152
rect 33066 33216 33382 33217
rect 33066 33152 33072 33216
rect 33136 33152 33152 33216
rect 33216 33152 33232 33216
rect 33296 33152 33312 33216
rect 33376 33152 33382 33216
rect 33066 33151 33382 33152
rect 3006 32672 3322 32673
rect 3006 32608 3012 32672
rect 3076 32608 3092 32672
rect 3156 32608 3172 32672
rect 3236 32608 3252 32672
rect 3316 32608 3322 32672
rect 3006 32607 3322 32608
rect 33726 32672 34042 32673
rect 33726 32608 33732 32672
rect 33796 32608 33812 32672
rect 33876 32608 33892 32672
rect 33956 32608 33972 32672
rect 34036 32608 34042 32672
rect 33726 32607 34042 32608
rect 2346 32128 2662 32129
rect 2346 32064 2352 32128
rect 2416 32064 2432 32128
rect 2496 32064 2512 32128
rect 2576 32064 2592 32128
rect 2656 32064 2662 32128
rect 2346 32063 2662 32064
rect 33066 32128 33382 32129
rect 33066 32064 33072 32128
rect 33136 32064 33152 32128
rect 33216 32064 33232 32128
rect 33296 32064 33312 32128
rect 33376 32064 33382 32128
rect 33066 32063 33382 32064
rect 3006 31584 3322 31585
rect 3006 31520 3012 31584
rect 3076 31520 3092 31584
rect 3156 31520 3172 31584
rect 3236 31520 3252 31584
rect 3316 31520 3322 31584
rect 3006 31519 3322 31520
rect 33726 31584 34042 31585
rect 33726 31520 33732 31584
rect 33796 31520 33812 31584
rect 33876 31520 33892 31584
rect 33956 31520 33972 31584
rect 34036 31520 34042 31584
rect 33726 31519 34042 31520
rect 2346 31040 2662 31041
rect 2346 30976 2352 31040
rect 2416 30976 2432 31040
rect 2496 30976 2512 31040
rect 2576 30976 2592 31040
rect 2656 30976 2662 31040
rect 2346 30975 2662 30976
rect 33066 31040 33382 31041
rect 33066 30976 33072 31040
rect 33136 30976 33152 31040
rect 33216 30976 33232 31040
rect 33296 30976 33312 31040
rect 33376 30976 33382 31040
rect 33066 30975 33382 30976
rect 3006 30496 3322 30497
rect 3006 30432 3012 30496
rect 3076 30432 3092 30496
rect 3156 30432 3172 30496
rect 3236 30432 3252 30496
rect 3316 30432 3322 30496
rect 3006 30431 3322 30432
rect 33726 30496 34042 30497
rect 33726 30432 33732 30496
rect 33796 30432 33812 30496
rect 33876 30432 33892 30496
rect 33956 30432 33972 30496
rect 34036 30432 34042 30496
rect 33726 30431 34042 30432
rect 2346 29952 2662 29953
rect 2346 29888 2352 29952
rect 2416 29888 2432 29952
rect 2496 29888 2512 29952
rect 2576 29888 2592 29952
rect 2656 29888 2662 29952
rect 2346 29887 2662 29888
rect 33066 29952 33382 29953
rect 33066 29888 33072 29952
rect 33136 29888 33152 29952
rect 33216 29888 33232 29952
rect 33296 29888 33312 29952
rect 33376 29888 33382 29952
rect 33066 29887 33382 29888
rect 3006 29408 3322 29409
rect 3006 29344 3012 29408
rect 3076 29344 3092 29408
rect 3156 29344 3172 29408
rect 3236 29344 3252 29408
rect 3316 29344 3322 29408
rect 3006 29343 3322 29344
rect 33726 29408 34042 29409
rect 33726 29344 33732 29408
rect 33796 29344 33812 29408
rect 33876 29344 33892 29408
rect 33956 29344 33972 29408
rect 34036 29344 34042 29408
rect 33726 29343 34042 29344
rect 2346 28864 2662 28865
rect 2346 28800 2352 28864
rect 2416 28800 2432 28864
rect 2496 28800 2512 28864
rect 2576 28800 2592 28864
rect 2656 28800 2662 28864
rect 2346 28799 2662 28800
rect 33066 28864 33382 28865
rect 33066 28800 33072 28864
rect 33136 28800 33152 28864
rect 33216 28800 33232 28864
rect 33296 28800 33312 28864
rect 33376 28800 33382 28864
rect 33066 28799 33382 28800
rect 3006 28320 3322 28321
rect 3006 28256 3012 28320
rect 3076 28256 3092 28320
rect 3156 28256 3172 28320
rect 3236 28256 3252 28320
rect 3316 28256 3322 28320
rect 3006 28255 3322 28256
rect 33726 28320 34042 28321
rect 33726 28256 33732 28320
rect 33796 28256 33812 28320
rect 33876 28256 33892 28320
rect 33956 28256 33972 28320
rect 34036 28256 34042 28320
rect 33726 28255 34042 28256
rect 2346 27776 2662 27777
rect 2346 27712 2352 27776
rect 2416 27712 2432 27776
rect 2496 27712 2512 27776
rect 2576 27712 2592 27776
rect 2656 27712 2662 27776
rect 2346 27711 2662 27712
rect 33066 27776 33382 27777
rect 33066 27712 33072 27776
rect 33136 27712 33152 27776
rect 33216 27712 33232 27776
rect 33296 27712 33312 27776
rect 33376 27712 33382 27776
rect 33066 27711 33382 27712
rect 3006 27232 3322 27233
rect 3006 27168 3012 27232
rect 3076 27168 3092 27232
rect 3156 27168 3172 27232
rect 3236 27168 3252 27232
rect 3316 27168 3322 27232
rect 3006 27167 3322 27168
rect 33726 27232 34042 27233
rect 33726 27168 33732 27232
rect 33796 27168 33812 27232
rect 33876 27168 33892 27232
rect 33956 27168 33972 27232
rect 34036 27168 34042 27232
rect 33726 27167 34042 27168
rect 2346 26688 2662 26689
rect 2346 26624 2352 26688
rect 2416 26624 2432 26688
rect 2496 26624 2512 26688
rect 2576 26624 2592 26688
rect 2656 26624 2662 26688
rect 2346 26623 2662 26624
rect 33066 26688 33382 26689
rect 33066 26624 33072 26688
rect 33136 26624 33152 26688
rect 33216 26624 33232 26688
rect 33296 26624 33312 26688
rect 33376 26624 33382 26688
rect 33066 26623 33382 26624
rect 3006 26144 3322 26145
rect 3006 26080 3012 26144
rect 3076 26080 3092 26144
rect 3156 26080 3172 26144
rect 3236 26080 3252 26144
rect 3316 26080 3322 26144
rect 3006 26079 3322 26080
rect 33726 26144 34042 26145
rect 33726 26080 33732 26144
rect 33796 26080 33812 26144
rect 33876 26080 33892 26144
rect 33956 26080 33972 26144
rect 34036 26080 34042 26144
rect 33726 26079 34042 26080
rect 2346 25600 2662 25601
rect 2346 25536 2352 25600
rect 2416 25536 2432 25600
rect 2496 25536 2512 25600
rect 2576 25536 2592 25600
rect 2656 25536 2662 25600
rect 2346 25535 2662 25536
rect 33066 25600 33382 25601
rect 33066 25536 33072 25600
rect 33136 25536 33152 25600
rect 33216 25536 33232 25600
rect 33296 25536 33312 25600
rect 33376 25536 33382 25600
rect 33066 25535 33382 25536
rect 3006 25056 3322 25057
rect 3006 24992 3012 25056
rect 3076 24992 3092 25056
rect 3156 24992 3172 25056
rect 3236 24992 3252 25056
rect 3316 24992 3322 25056
rect 3006 24991 3322 24992
rect 33726 25056 34042 25057
rect 33726 24992 33732 25056
rect 33796 24992 33812 25056
rect 33876 24992 33892 25056
rect 33956 24992 33972 25056
rect 34036 24992 34042 25056
rect 33726 24991 34042 24992
rect 2346 24512 2662 24513
rect 2346 24448 2352 24512
rect 2416 24448 2432 24512
rect 2496 24448 2512 24512
rect 2576 24448 2592 24512
rect 2656 24448 2662 24512
rect 2346 24447 2662 24448
rect 33066 24512 33382 24513
rect 33066 24448 33072 24512
rect 33136 24448 33152 24512
rect 33216 24448 33232 24512
rect 33296 24448 33312 24512
rect 33376 24448 33382 24512
rect 33066 24447 33382 24448
rect 3006 23968 3322 23969
rect 3006 23904 3012 23968
rect 3076 23904 3092 23968
rect 3156 23904 3172 23968
rect 3236 23904 3252 23968
rect 3316 23904 3322 23968
rect 3006 23903 3322 23904
rect 33726 23968 34042 23969
rect 33726 23904 33732 23968
rect 33796 23904 33812 23968
rect 33876 23904 33892 23968
rect 33956 23904 33972 23968
rect 34036 23904 34042 23968
rect 33726 23903 34042 23904
rect 2346 23424 2662 23425
rect 2346 23360 2352 23424
rect 2416 23360 2432 23424
rect 2496 23360 2512 23424
rect 2576 23360 2592 23424
rect 2656 23360 2662 23424
rect 2346 23359 2662 23360
rect 33066 23424 33382 23425
rect 33066 23360 33072 23424
rect 33136 23360 33152 23424
rect 33216 23360 33232 23424
rect 33296 23360 33312 23424
rect 33376 23360 33382 23424
rect 33066 23359 33382 23360
rect 3006 22880 3322 22881
rect 3006 22816 3012 22880
rect 3076 22816 3092 22880
rect 3156 22816 3172 22880
rect 3236 22816 3252 22880
rect 3316 22816 3322 22880
rect 3006 22815 3322 22816
rect 33726 22880 34042 22881
rect 33726 22816 33732 22880
rect 33796 22816 33812 22880
rect 33876 22816 33892 22880
rect 33956 22816 33972 22880
rect 34036 22816 34042 22880
rect 33726 22815 34042 22816
rect 2346 22336 2662 22337
rect 2346 22272 2352 22336
rect 2416 22272 2432 22336
rect 2496 22272 2512 22336
rect 2576 22272 2592 22336
rect 2656 22272 2662 22336
rect 2346 22271 2662 22272
rect 33066 22336 33382 22337
rect 33066 22272 33072 22336
rect 33136 22272 33152 22336
rect 33216 22272 33232 22336
rect 33296 22272 33312 22336
rect 33376 22272 33382 22336
rect 33066 22271 33382 22272
rect 3006 21792 3322 21793
rect 3006 21728 3012 21792
rect 3076 21728 3092 21792
rect 3156 21728 3172 21792
rect 3236 21728 3252 21792
rect 3316 21728 3322 21792
rect 3006 21727 3322 21728
rect 33726 21792 34042 21793
rect 33726 21728 33732 21792
rect 33796 21728 33812 21792
rect 33876 21728 33892 21792
rect 33956 21728 33972 21792
rect 34036 21728 34042 21792
rect 33726 21727 34042 21728
rect 2346 21248 2662 21249
rect 2346 21184 2352 21248
rect 2416 21184 2432 21248
rect 2496 21184 2512 21248
rect 2576 21184 2592 21248
rect 2656 21184 2662 21248
rect 2346 21183 2662 21184
rect 33066 21248 33382 21249
rect 33066 21184 33072 21248
rect 33136 21184 33152 21248
rect 33216 21184 33232 21248
rect 33296 21184 33312 21248
rect 33376 21184 33382 21248
rect 33066 21183 33382 21184
rect 3006 20704 3322 20705
rect 3006 20640 3012 20704
rect 3076 20640 3092 20704
rect 3156 20640 3172 20704
rect 3236 20640 3252 20704
rect 3316 20640 3322 20704
rect 3006 20639 3322 20640
rect 33726 20704 34042 20705
rect 33726 20640 33732 20704
rect 33796 20640 33812 20704
rect 33876 20640 33892 20704
rect 33956 20640 33972 20704
rect 34036 20640 34042 20704
rect 33726 20639 34042 20640
rect 2346 20160 2662 20161
rect 2346 20096 2352 20160
rect 2416 20096 2432 20160
rect 2496 20096 2512 20160
rect 2576 20096 2592 20160
rect 2656 20096 2662 20160
rect 2346 20095 2662 20096
rect 33066 20160 33382 20161
rect 33066 20096 33072 20160
rect 33136 20096 33152 20160
rect 33216 20096 33232 20160
rect 33296 20096 33312 20160
rect 33376 20096 33382 20160
rect 33066 20095 33382 20096
rect 3006 19616 3322 19617
rect 3006 19552 3012 19616
rect 3076 19552 3092 19616
rect 3156 19552 3172 19616
rect 3236 19552 3252 19616
rect 3316 19552 3322 19616
rect 3006 19551 3322 19552
rect 33726 19616 34042 19617
rect 33726 19552 33732 19616
rect 33796 19552 33812 19616
rect 33876 19552 33892 19616
rect 33956 19552 33972 19616
rect 34036 19552 34042 19616
rect 33726 19551 34042 19552
rect 2346 19072 2662 19073
rect 2346 19008 2352 19072
rect 2416 19008 2432 19072
rect 2496 19008 2512 19072
rect 2576 19008 2592 19072
rect 2656 19008 2662 19072
rect 2346 19007 2662 19008
rect 33066 19072 33382 19073
rect 33066 19008 33072 19072
rect 33136 19008 33152 19072
rect 33216 19008 33232 19072
rect 33296 19008 33312 19072
rect 33376 19008 33382 19072
rect 33066 19007 33382 19008
rect 3006 18528 3322 18529
rect 3006 18464 3012 18528
rect 3076 18464 3092 18528
rect 3156 18464 3172 18528
rect 3236 18464 3252 18528
rect 3316 18464 3322 18528
rect 3006 18463 3322 18464
rect 33726 18528 34042 18529
rect 33726 18464 33732 18528
rect 33796 18464 33812 18528
rect 33876 18464 33892 18528
rect 33956 18464 33972 18528
rect 34036 18464 34042 18528
rect 33726 18463 34042 18464
rect 2346 17984 2662 17985
rect 2346 17920 2352 17984
rect 2416 17920 2432 17984
rect 2496 17920 2512 17984
rect 2576 17920 2592 17984
rect 2656 17920 2662 17984
rect 2346 17919 2662 17920
rect 33066 17984 33382 17985
rect 33066 17920 33072 17984
rect 33136 17920 33152 17984
rect 33216 17920 33232 17984
rect 33296 17920 33312 17984
rect 33376 17920 33382 17984
rect 33066 17919 33382 17920
rect 3006 17440 3322 17441
rect 3006 17376 3012 17440
rect 3076 17376 3092 17440
rect 3156 17376 3172 17440
rect 3236 17376 3252 17440
rect 3316 17376 3322 17440
rect 3006 17375 3322 17376
rect 33726 17440 34042 17441
rect 33726 17376 33732 17440
rect 33796 17376 33812 17440
rect 33876 17376 33892 17440
rect 33956 17376 33972 17440
rect 34036 17376 34042 17440
rect 33726 17375 34042 17376
rect 2346 16896 2662 16897
rect 2346 16832 2352 16896
rect 2416 16832 2432 16896
rect 2496 16832 2512 16896
rect 2576 16832 2592 16896
rect 2656 16832 2662 16896
rect 2346 16831 2662 16832
rect 33066 16896 33382 16897
rect 33066 16832 33072 16896
rect 33136 16832 33152 16896
rect 33216 16832 33232 16896
rect 33296 16832 33312 16896
rect 33376 16832 33382 16896
rect 33066 16831 33382 16832
rect 3006 16352 3322 16353
rect 3006 16288 3012 16352
rect 3076 16288 3092 16352
rect 3156 16288 3172 16352
rect 3236 16288 3252 16352
rect 3316 16288 3322 16352
rect 3006 16287 3322 16288
rect 33726 16352 34042 16353
rect 33726 16288 33732 16352
rect 33796 16288 33812 16352
rect 33876 16288 33892 16352
rect 33956 16288 33972 16352
rect 34036 16288 34042 16352
rect 33726 16287 34042 16288
rect 2346 15808 2662 15809
rect 2346 15744 2352 15808
rect 2416 15744 2432 15808
rect 2496 15744 2512 15808
rect 2576 15744 2592 15808
rect 2656 15744 2662 15808
rect 2346 15743 2662 15744
rect 33066 15808 33382 15809
rect 33066 15744 33072 15808
rect 33136 15744 33152 15808
rect 33216 15744 33232 15808
rect 33296 15744 33312 15808
rect 33376 15744 33382 15808
rect 33066 15743 33382 15744
rect 3006 15264 3322 15265
rect 3006 15200 3012 15264
rect 3076 15200 3092 15264
rect 3156 15200 3172 15264
rect 3236 15200 3252 15264
rect 3316 15200 3322 15264
rect 3006 15199 3322 15200
rect 33726 15264 34042 15265
rect 33726 15200 33732 15264
rect 33796 15200 33812 15264
rect 33876 15200 33892 15264
rect 33956 15200 33972 15264
rect 34036 15200 34042 15264
rect 33726 15199 34042 15200
rect 56501 15058 56567 15061
rect 59200 15058 60000 15088
rect 56501 15056 60000 15058
rect 56501 15000 56506 15056
rect 56562 15000 60000 15056
rect 56501 14998 60000 15000
rect 56501 14995 56567 14998
rect 59200 14968 60000 14998
rect 2346 14720 2662 14721
rect 2346 14656 2352 14720
rect 2416 14656 2432 14720
rect 2496 14656 2512 14720
rect 2576 14656 2592 14720
rect 2656 14656 2662 14720
rect 2346 14655 2662 14656
rect 33066 14720 33382 14721
rect 33066 14656 33072 14720
rect 33136 14656 33152 14720
rect 33216 14656 33232 14720
rect 33296 14656 33312 14720
rect 33376 14656 33382 14720
rect 33066 14655 33382 14656
rect 3006 14176 3322 14177
rect 3006 14112 3012 14176
rect 3076 14112 3092 14176
rect 3156 14112 3172 14176
rect 3236 14112 3252 14176
rect 3316 14112 3322 14176
rect 3006 14111 3322 14112
rect 33726 14176 34042 14177
rect 33726 14112 33732 14176
rect 33796 14112 33812 14176
rect 33876 14112 33892 14176
rect 33956 14112 33972 14176
rect 34036 14112 34042 14176
rect 33726 14111 34042 14112
rect 2346 13632 2662 13633
rect 2346 13568 2352 13632
rect 2416 13568 2432 13632
rect 2496 13568 2512 13632
rect 2576 13568 2592 13632
rect 2656 13568 2662 13632
rect 2346 13567 2662 13568
rect 33066 13632 33382 13633
rect 33066 13568 33072 13632
rect 33136 13568 33152 13632
rect 33216 13568 33232 13632
rect 33296 13568 33312 13632
rect 33376 13568 33382 13632
rect 33066 13567 33382 13568
rect 3006 13088 3322 13089
rect 3006 13024 3012 13088
rect 3076 13024 3092 13088
rect 3156 13024 3172 13088
rect 3236 13024 3252 13088
rect 3316 13024 3322 13088
rect 3006 13023 3322 13024
rect 33726 13088 34042 13089
rect 33726 13024 33732 13088
rect 33796 13024 33812 13088
rect 33876 13024 33892 13088
rect 33956 13024 33972 13088
rect 34036 13024 34042 13088
rect 33726 13023 34042 13024
rect 2346 12544 2662 12545
rect 2346 12480 2352 12544
rect 2416 12480 2432 12544
rect 2496 12480 2512 12544
rect 2576 12480 2592 12544
rect 2656 12480 2662 12544
rect 2346 12479 2662 12480
rect 33066 12544 33382 12545
rect 33066 12480 33072 12544
rect 33136 12480 33152 12544
rect 33216 12480 33232 12544
rect 33296 12480 33312 12544
rect 33376 12480 33382 12544
rect 33066 12479 33382 12480
rect 3006 12000 3322 12001
rect 3006 11936 3012 12000
rect 3076 11936 3092 12000
rect 3156 11936 3172 12000
rect 3236 11936 3252 12000
rect 3316 11936 3322 12000
rect 3006 11935 3322 11936
rect 33726 12000 34042 12001
rect 33726 11936 33732 12000
rect 33796 11936 33812 12000
rect 33876 11936 33892 12000
rect 33956 11936 33972 12000
rect 34036 11936 34042 12000
rect 33726 11935 34042 11936
rect 2346 11456 2662 11457
rect 2346 11392 2352 11456
rect 2416 11392 2432 11456
rect 2496 11392 2512 11456
rect 2576 11392 2592 11456
rect 2656 11392 2662 11456
rect 2346 11391 2662 11392
rect 33066 11456 33382 11457
rect 33066 11392 33072 11456
rect 33136 11392 33152 11456
rect 33216 11392 33232 11456
rect 33296 11392 33312 11456
rect 33376 11392 33382 11456
rect 33066 11391 33382 11392
rect 3006 10912 3322 10913
rect 3006 10848 3012 10912
rect 3076 10848 3092 10912
rect 3156 10848 3172 10912
rect 3236 10848 3252 10912
rect 3316 10848 3322 10912
rect 3006 10847 3322 10848
rect 33726 10912 34042 10913
rect 33726 10848 33732 10912
rect 33796 10848 33812 10912
rect 33876 10848 33892 10912
rect 33956 10848 33972 10912
rect 34036 10848 34042 10912
rect 33726 10847 34042 10848
rect 2346 10368 2662 10369
rect 2346 10304 2352 10368
rect 2416 10304 2432 10368
rect 2496 10304 2512 10368
rect 2576 10304 2592 10368
rect 2656 10304 2662 10368
rect 2346 10303 2662 10304
rect 33066 10368 33382 10369
rect 33066 10304 33072 10368
rect 33136 10304 33152 10368
rect 33216 10304 33232 10368
rect 33296 10304 33312 10368
rect 33376 10304 33382 10368
rect 33066 10303 33382 10304
rect 3006 9824 3322 9825
rect 3006 9760 3012 9824
rect 3076 9760 3092 9824
rect 3156 9760 3172 9824
rect 3236 9760 3252 9824
rect 3316 9760 3322 9824
rect 3006 9759 3322 9760
rect 33726 9824 34042 9825
rect 33726 9760 33732 9824
rect 33796 9760 33812 9824
rect 33876 9760 33892 9824
rect 33956 9760 33972 9824
rect 34036 9760 34042 9824
rect 33726 9759 34042 9760
rect 2346 9280 2662 9281
rect 2346 9216 2352 9280
rect 2416 9216 2432 9280
rect 2496 9216 2512 9280
rect 2576 9216 2592 9280
rect 2656 9216 2662 9280
rect 2346 9215 2662 9216
rect 33066 9280 33382 9281
rect 33066 9216 33072 9280
rect 33136 9216 33152 9280
rect 33216 9216 33232 9280
rect 33296 9216 33312 9280
rect 33376 9216 33382 9280
rect 33066 9215 33382 9216
rect 3006 8736 3322 8737
rect 3006 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3322 8736
rect 3006 8671 3322 8672
rect 33726 8736 34042 8737
rect 33726 8672 33732 8736
rect 33796 8672 33812 8736
rect 33876 8672 33892 8736
rect 33956 8672 33972 8736
rect 34036 8672 34042 8736
rect 33726 8671 34042 8672
rect 2346 8192 2662 8193
rect 2346 8128 2352 8192
rect 2416 8128 2432 8192
rect 2496 8128 2512 8192
rect 2576 8128 2592 8192
rect 2656 8128 2662 8192
rect 2346 8127 2662 8128
rect 33066 8192 33382 8193
rect 33066 8128 33072 8192
rect 33136 8128 33152 8192
rect 33216 8128 33232 8192
rect 33296 8128 33312 8192
rect 33376 8128 33382 8192
rect 33066 8127 33382 8128
rect 3006 7648 3322 7649
rect 3006 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3322 7648
rect 3006 7583 3322 7584
rect 33726 7648 34042 7649
rect 33726 7584 33732 7648
rect 33796 7584 33812 7648
rect 33876 7584 33892 7648
rect 33956 7584 33972 7648
rect 34036 7584 34042 7648
rect 33726 7583 34042 7584
rect 2346 7104 2662 7105
rect 2346 7040 2352 7104
rect 2416 7040 2432 7104
rect 2496 7040 2512 7104
rect 2576 7040 2592 7104
rect 2656 7040 2662 7104
rect 2346 7039 2662 7040
rect 33066 7104 33382 7105
rect 33066 7040 33072 7104
rect 33136 7040 33152 7104
rect 33216 7040 33232 7104
rect 33296 7040 33312 7104
rect 33376 7040 33382 7104
rect 33066 7039 33382 7040
rect 3006 6560 3322 6561
rect 3006 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3322 6560
rect 3006 6495 3322 6496
rect 33726 6560 34042 6561
rect 33726 6496 33732 6560
rect 33796 6496 33812 6560
rect 33876 6496 33892 6560
rect 33956 6496 33972 6560
rect 34036 6496 34042 6560
rect 33726 6495 34042 6496
rect 2346 6016 2662 6017
rect 2346 5952 2352 6016
rect 2416 5952 2432 6016
rect 2496 5952 2512 6016
rect 2576 5952 2592 6016
rect 2656 5952 2662 6016
rect 2346 5951 2662 5952
rect 33066 6016 33382 6017
rect 33066 5952 33072 6016
rect 33136 5952 33152 6016
rect 33216 5952 33232 6016
rect 33296 5952 33312 6016
rect 33376 5952 33382 6016
rect 33066 5951 33382 5952
rect 3006 5472 3322 5473
rect 3006 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3322 5472
rect 3006 5407 3322 5408
rect 33726 5472 34042 5473
rect 33726 5408 33732 5472
rect 33796 5408 33812 5472
rect 33876 5408 33892 5472
rect 33956 5408 33972 5472
rect 34036 5408 34042 5472
rect 33726 5407 34042 5408
rect 2346 4928 2662 4929
rect 2346 4864 2352 4928
rect 2416 4864 2432 4928
rect 2496 4864 2512 4928
rect 2576 4864 2592 4928
rect 2656 4864 2662 4928
rect 2346 4863 2662 4864
rect 33066 4928 33382 4929
rect 33066 4864 33072 4928
rect 33136 4864 33152 4928
rect 33216 4864 33232 4928
rect 33296 4864 33312 4928
rect 33376 4864 33382 4928
rect 33066 4863 33382 4864
rect 3006 4384 3322 4385
rect 3006 4320 3012 4384
rect 3076 4320 3092 4384
rect 3156 4320 3172 4384
rect 3236 4320 3252 4384
rect 3316 4320 3322 4384
rect 3006 4319 3322 4320
rect 33726 4384 34042 4385
rect 33726 4320 33732 4384
rect 33796 4320 33812 4384
rect 33876 4320 33892 4384
rect 33956 4320 33972 4384
rect 34036 4320 34042 4384
rect 33726 4319 34042 4320
rect 2346 3840 2662 3841
rect 2346 3776 2352 3840
rect 2416 3776 2432 3840
rect 2496 3776 2512 3840
rect 2576 3776 2592 3840
rect 2656 3776 2662 3840
rect 2346 3775 2662 3776
rect 33066 3840 33382 3841
rect 33066 3776 33072 3840
rect 33136 3776 33152 3840
rect 33216 3776 33232 3840
rect 33296 3776 33312 3840
rect 33376 3776 33382 3840
rect 33066 3775 33382 3776
rect 3006 3296 3322 3297
rect 3006 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3322 3296
rect 3006 3231 3322 3232
rect 33726 3296 34042 3297
rect 33726 3232 33732 3296
rect 33796 3232 33812 3296
rect 33876 3232 33892 3296
rect 33956 3232 33972 3296
rect 34036 3232 34042 3296
rect 33726 3231 34042 3232
rect 2346 2752 2662 2753
rect 2346 2688 2352 2752
rect 2416 2688 2432 2752
rect 2496 2688 2512 2752
rect 2576 2688 2592 2752
rect 2656 2688 2662 2752
rect 2346 2687 2662 2688
rect 33066 2752 33382 2753
rect 33066 2688 33072 2752
rect 33136 2688 33152 2752
rect 33216 2688 33232 2752
rect 33296 2688 33312 2752
rect 33376 2688 33382 2752
rect 33066 2687 33382 2688
rect 3006 2208 3322 2209
rect 3006 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3322 2208
rect 3006 2143 3322 2144
rect 33726 2208 34042 2209
rect 33726 2144 33732 2208
rect 33796 2144 33812 2208
rect 33876 2144 33892 2208
rect 33956 2144 33972 2208
rect 34036 2144 34042 2208
rect 33726 2143 34042 2144
<< via3 >>
rect 3012 57692 3076 57696
rect 3012 57636 3016 57692
rect 3016 57636 3072 57692
rect 3072 57636 3076 57692
rect 3012 57632 3076 57636
rect 3092 57692 3156 57696
rect 3092 57636 3096 57692
rect 3096 57636 3152 57692
rect 3152 57636 3156 57692
rect 3092 57632 3156 57636
rect 3172 57692 3236 57696
rect 3172 57636 3176 57692
rect 3176 57636 3232 57692
rect 3232 57636 3236 57692
rect 3172 57632 3236 57636
rect 3252 57692 3316 57696
rect 3252 57636 3256 57692
rect 3256 57636 3312 57692
rect 3312 57636 3316 57692
rect 3252 57632 3316 57636
rect 33732 57692 33796 57696
rect 33732 57636 33736 57692
rect 33736 57636 33792 57692
rect 33792 57636 33796 57692
rect 33732 57632 33796 57636
rect 33812 57692 33876 57696
rect 33812 57636 33816 57692
rect 33816 57636 33872 57692
rect 33872 57636 33876 57692
rect 33812 57632 33876 57636
rect 33892 57692 33956 57696
rect 33892 57636 33896 57692
rect 33896 57636 33952 57692
rect 33952 57636 33956 57692
rect 33892 57632 33956 57636
rect 33972 57692 34036 57696
rect 33972 57636 33976 57692
rect 33976 57636 34032 57692
rect 34032 57636 34036 57692
rect 33972 57632 34036 57636
rect 2352 57148 2416 57152
rect 2352 57092 2356 57148
rect 2356 57092 2412 57148
rect 2412 57092 2416 57148
rect 2352 57088 2416 57092
rect 2432 57148 2496 57152
rect 2432 57092 2436 57148
rect 2436 57092 2492 57148
rect 2492 57092 2496 57148
rect 2432 57088 2496 57092
rect 2512 57148 2576 57152
rect 2512 57092 2516 57148
rect 2516 57092 2572 57148
rect 2572 57092 2576 57148
rect 2512 57088 2576 57092
rect 2592 57148 2656 57152
rect 2592 57092 2596 57148
rect 2596 57092 2652 57148
rect 2652 57092 2656 57148
rect 2592 57088 2656 57092
rect 33072 57148 33136 57152
rect 33072 57092 33076 57148
rect 33076 57092 33132 57148
rect 33132 57092 33136 57148
rect 33072 57088 33136 57092
rect 33152 57148 33216 57152
rect 33152 57092 33156 57148
rect 33156 57092 33212 57148
rect 33212 57092 33216 57148
rect 33152 57088 33216 57092
rect 33232 57148 33296 57152
rect 33232 57092 33236 57148
rect 33236 57092 33292 57148
rect 33292 57092 33296 57148
rect 33232 57088 33296 57092
rect 33312 57148 33376 57152
rect 33312 57092 33316 57148
rect 33316 57092 33372 57148
rect 33372 57092 33376 57148
rect 33312 57088 33376 57092
rect 3012 56604 3076 56608
rect 3012 56548 3016 56604
rect 3016 56548 3072 56604
rect 3072 56548 3076 56604
rect 3012 56544 3076 56548
rect 3092 56604 3156 56608
rect 3092 56548 3096 56604
rect 3096 56548 3152 56604
rect 3152 56548 3156 56604
rect 3092 56544 3156 56548
rect 3172 56604 3236 56608
rect 3172 56548 3176 56604
rect 3176 56548 3232 56604
rect 3232 56548 3236 56604
rect 3172 56544 3236 56548
rect 3252 56604 3316 56608
rect 3252 56548 3256 56604
rect 3256 56548 3312 56604
rect 3312 56548 3316 56604
rect 3252 56544 3316 56548
rect 33732 56604 33796 56608
rect 33732 56548 33736 56604
rect 33736 56548 33792 56604
rect 33792 56548 33796 56604
rect 33732 56544 33796 56548
rect 33812 56604 33876 56608
rect 33812 56548 33816 56604
rect 33816 56548 33872 56604
rect 33872 56548 33876 56604
rect 33812 56544 33876 56548
rect 33892 56604 33956 56608
rect 33892 56548 33896 56604
rect 33896 56548 33952 56604
rect 33952 56548 33956 56604
rect 33892 56544 33956 56548
rect 33972 56604 34036 56608
rect 33972 56548 33976 56604
rect 33976 56548 34032 56604
rect 34032 56548 34036 56604
rect 33972 56544 34036 56548
rect 2352 56060 2416 56064
rect 2352 56004 2356 56060
rect 2356 56004 2412 56060
rect 2412 56004 2416 56060
rect 2352 56000 2416 56004
rect 2432 56060 2496 56064
rect 2432 56004 2436 56060
rect 2436 56004 2492 56060
rect 2492 56004 2496 56060
rect 2432 56000 2496 56004
rect 2512 56060 2576 56064
rect 2512 56004 2516 56060
rect 2516 56004 2572 56060
rect 2572 56004 2576 56060
rect 2512 56000 2576 56004
rect 2592 56060 2656 56064
rect 2592 56004 2596 56060
rect 2596 56004 2652 56060
rect 2652 56004 2656 56060
rect 2592 56000 2656 56004
rect 33072 56060 33136 56064
rect 33072 56004 33076 56060
rect 33076 56004 33132 56060
rect 33132 56004 33136 56060
rect 33072 56000 33136 56004
rect 33152 56060 33216 56064
rect 33152 56004 33156 56060
rect 33156 56004 33212 56060
rect 33212 56004 33216 56060
rect 33152 56000 33216 56004
rect 33232 56060 33296 56064
rect 33232 56004 33236 56060
rect 33236 56004 33292 56060
rect 33292 56004 33296 56060
rect 33232 56000 33296 56004
rect 33312 56060 33376 56064
rect 33312 56004 33316 56060
rect 33316 56004 33372 56060
rect 33372 56004 33376 56060
rect 33312 56000 33376 56004
rect 3012 55516 3076 55520
rect 3012 55460 3016 55516
rect 3016 55460 3072 55516
rect 3072 55460 3076 55516
rect 3012 55456 3076 55460
rect 3092 55516 3156 55520
rect 3092 55460 3096 55516
rect 3096 55460 3152 55516
rect 3152 55460 3156 55516
rect 3092 55456 3156 55460
rect 3172 55516 3236 55520
rect 3172 55460 3176 55516
rect 3176 55460 3232 55516
rect 3232 55460 3236 55516
rect 3172 55456 3236 55460
rect 3252 55516 3316 55520
rect 3252 55460 3256 55516
rect 3256 55460 3312 55516
rect 3312 55460 3316 55516
rect 3252 55456 3316 55460
rect 33732 55516 33796 55520
rect 33732 55460 33736 55516
rect 33736 55460 33792 55516
rect 33792 55460 33796 55516
rect 33732 55456 33796 55460
rect 33812 55516 33876 55520
rect 33812 55460 33816 55516
rect 33816 55460 33872 55516
rect 33872 55460 33876 55516
rect 33812 55456 33876 55460
rect 33892 55516 33956 55520
rect 33892 55460 33896 55516
rect 33896 55460 33952 55516
rect 33952 55460 33956 55516
rect 33892 55456 33956 55460
rect 33972 55516 34036 55520
rect 33972 55460 33976 55516
rect 33976 55460 34032 55516
rect 34032 55460 34036 55516
rect 33972 55456 34036 55460
rect 2352 54972 2416 54976
rect 2352 54916 2356 54972
rect 2356 54916 2412 54972
rect 2412 54916 2416 54972
rect 2352 54912 2416 54916
rect 2432 54972 2496 54976
rect 2432 54916 2436 54972
rect 2436 54916 2492 54972
rect 2492 54916 2496 54972
rect 2432 54912 2496 54916
rect 2512 54972 2576 54976
rect 2512 54916 2516 54972
rect 2516 54916 2572 54972
rect 2572 54916 2576 54972
rect 2512 54912 2576 54916
rect 2592 54972 2656 54976
rect 2592 54916 2596 54972
rect 2596 54916 2652 54972
rect 2652 54916 2656 54972
rect 2592 54912 2656 54916
rect 33072 54972 33136 54976
rect 33072 54916 33076 54972
rect 33076 54916 33132 54972
rect 33132 54916 33136 54972
rect 33072 54912 33136 54916
rect 33152 54972 33216 54976
rect 33152 54916 33156 54972
rect 33156 54916 33212 54972
rect 33212 54916 33216 54972
rect 33152 54912 33216 54916
rect 33232 54972 33296 54976
rect 33232 54916 33236 54972
rect 33236 54916 33292 54972
rect 33292 54916 33296 54972
rect 33232 54912 33296 54916
rect 33312 54972 33376 54976
rect 33312 54916 33316 54972
rect 33316 54916 33372 54972
rect 33372 54916 33376 54972
rect 33312 54912 33376 54916
rect 3012 54428 3076 54432
rect 3012 54372 3016 54428
rect 3016 54372 3072 54428
rect 3072 54372 3076 54428
rect 3012 54368 3076 54372
rect 3092 54428 3156 54432
rect 3092 54372 3096 54428
rect 3096 54372 3152 54428
rect 3152 54372 3156 54428
rect 3092 54368 3156 54372
rect 3172 54428 3236 54432
rect 3172 54372 3176 54428
rect 3176 54372 3232 54428
rect 3232 54372 3236 54428
rect 3172 54368 3236 54372
rect 3252 54428 3316 54432
rect 3252 54372 3256 54428
rect 3256 54372 3312 54428
rect 3312 54372 3316 54428
rect 3252 54368 3316 54372
rect 33732 54428 33796 54432
rect 33732 54372 33736 54428
rect 33736 54372 33792 54428
rect 33792 54372 33796 54428
rect 33732 54368 33796 54372
rect 33812 54428 33876 54432
rect 33812 54372 33816 54428
rect 33816 54372 33872 54428
rect 33872 54372 33876 54428
rect 33812 54368 33876 54372
rect 33892 54428 33956 54432
rect 33892 54372 33896 54428
rect 33896 54372 33952 54428
rect 33952 54372 33956 54428
rect 33892 54368 33956 54372
rect 33972 54428 34036 54432
rect 33972 54372 33976 54428
rect 33976 54372 34032 54428
rect 34032 54372 34036 54428
rect 33972 54368 34036 54372
rect 2352 53884 2416 53888
rect 2352 53828 2356 53884
rect 2356 53828 2412 53884
rect 2412 53828 2416 53884
rect 2352 53824 2416 53828
rect 2432 53884 2496 53888
rect 2432 53828 2436 53884
rect 2436 53828 2492 53884
rect 2492 53828 2496 53884
rect 2432 53824 2496 53828
rect 2512 53884 2576 53888
rect 2512 53828 2516 53884
rect 2516 53828 2572 53884
rect 2572 53828 2576 53884
rect 2512 53824 2576 53828
rect 2592 53884 2656 53888
rect 2592 53828 2596 53884
rect 2596 53828 2652 53884
rect 2652 53828 2656 53884
rect 2592 53824 2656 53828
rect 33072 53884 33136 53888
rect 33072 53828 33076 53884
rect 33076 53828 33132 53884
rect 33132 53828 33136 53884
rect 33072 53824 33136 53828
rect 33152 53884 33216 53888
rect 33152 53828 33156 53884
rect 33156 53828 33212 53884
rect 33212 53828 33216 53884
rect 33152 53824 33216 53828
rect 33232 53884 33296 53888
rect 33232 53828 33236 53884
rect 33236 53828 33292 53884
rect 33292 53828 33296 53884
rect 33232 53824 33296 53828
rect 33312 53884 33376 53888
rect 33312 53828 33316 53884
rect 33316 53828 33372 53884
rect 33372 53828 33376 53884
rect 33312 53824 33376 53828
rect 3012 53340 3076 53344
rect 3012 53284 3016 53340
rect 3016 53284 3072 53340
rect 3072 53284 3076 53340
rect 3012 53280 3076 53284
rect 3092 53340 3156 53344
rect 3092 53284 3096 53340
rect 3096 53284 3152 53340
rect 3152 53284 3156 53340
rect 3092 53280 3156 53284
rect 3172 53340 3236 53344
rect 3172 53284 3176 53340
rect 3176 53284 3232 53340
rect 3232 53284 3236 53340
rect 3172 53280 3236 53284
rect 3252 53340 3316 53344
rect 3252 53284 3256 53340
rect 3256 53284 3312 53340
rect 3312 53284 3316 53340
rect 3252 53280 3316 53284
rect 33732 53340 33796 53344
rect 33732 53284 33736 53340
rect 33736 53284 33792 53340
rect 33792 53284 33796 53340
rect 33732 53280 33796 53284
rect 33812 53340 33876 53344
rect 33812 53284 33816 53340
rect 33816 53284 33872 53340
rect 33872 53284 33876 53340
rect 33812 53280 33876 53284
rect 33892 53340 33956 53344
rect 33892 53284 33896 53340
rect 33896 53284 33952 53340
rect 33952 53284 33956 53340
rect 33892 53280 33956 53284
rect 33972 53340 34036 53344
rect 33972 53284 33976 53340
rect 33976 53284 34032 53340
rect 34032 53284 34036 53340
rect 33972 53280 34036 53284
rect 2352 52796 2416 52800
rect 2352 52740 2356 52796
rect 2356 52740 2412 52796
rect 2412 52740 2416 52796
rect 2352 52736 2416 52740
rect 2432 52796 2496 52800
rect 2432 52740 2436 52796
rect 2436 52740 2492 52796
rect 2492 52740 2496 52796
rect 2432 52736 2496 52740
rect 2512 52796 2576 52800
rect 2512 52740 2516 52796
rect 2516 52740 2572 52796
rect 2572 52740 2576 52796
rect 2512 52736 2576 52740
rect 2592 52796 2656 52800
rect 2592 52740 2596 52796
rect 2596 52740 2652 52796
rect 2652 52740 2656 52796
rect 2592 52736 2656 52740
rect 33072 52796 33136 52800
rect 33072 52740 33076 52796
rect 33076 52740 33132 52796
rect 33132 52740 33136 52796
rect 33072 52736 33136 52740
rect 33152 52796 33216 52800
rect 33152 52740 33156 52796
rect 33156 52740 33212 52796
rect 33212 52740 33216 52796
rect 33152 52736 33216 52740
rect 33232 52796 33296 52800
rect 33232 52740 33236 52796
rect 33236 52740 33292 52796
rect 33292 52740 33296 52796
rect 33232 52736 33296 52740
rect 33312 52796 33376 52800
rect 33312 52740 33316 52796
rect 33316 52740 33372 52796
rect 33372 52740 33376 52796
rect 33312 52736 33376 52740
rect 3012 52252 3076 52256
rect 3012 52196 3016 52252
rect 3016 52196 3072 52252
rect 3072 52196 3076 52252
rect 3012 52192 3076 52196
rect 3092 52252 3156 52256
rect 3092 52196 3096 52252
rect 3096 52196 3152 52252
rect 3152 52196 3156 52252
rect 3092 52192 3156 52196
rect 3172 52252 3236 52256
rect 3172 52196 3176 52252
rect 3176 52196 3232 52252
rect 3232 52196 3236 52252
rect 3172 52192 3236 52196
rect 3252 52252 3316 52256
rect 3252 52196 3256 52252
rect 3256 52196 3312 52252
rect 3312 52196 3316 52252
rect 3252 52192 3316 52196
rect 33732 52252 33796 52256
rect 33732 52196 33736 52252
rect 33736 52196 33792 52252
rect 33792 52196 33796 52252
rect 33732 52192 33796 52196
rect 33812 52252 33876 52256
rect 33812 52196 33816 52252
rect 33816 52196 33872 52252
rect 33872 52196 33876 52252
rect 33812 52192 33876 52196
rect 33892 52252 33956 52256
rect 33892 52196 33896 52252
rect 33896 52196 33952 52252
rect 33952 52196 33956 52252
rect 33892 52192 33956 52196
rect 33972 52252 34036 52256
rect 33972 52196 33976 52252
rect 33976 52196 34032 52252
rect 34032 52196 34036 52252
rect 33972 52192 34036 52196
rect 2352 51708 2416 51712
rect 2352 51652 2356 51708
rect 2356 51652 2412 51708
rect 2412 51652 2416 51708
rect 2352 51648 2416 51652
rect 2432 51708 2496 51712
rect 2432 51652 2436 51708
rect 2436 51652 2492 51708
rect 2492 51652 2496 51708
rect 2432 51648 2496 51652
rect 2512 51708 2576 51712
rect 2512 51652 2516 51708
rect 2516 51652 2572 51708
rect 2572 51652 2576 51708
rect 2512 51648 2576 51652
rect 2592 51708 2656 51712
rect 2592 51652 2596 51708
rect 2596 51652 2652 51708
rect 2652 51652 2656 51708
rect 2592 51648 2656 51652
rect 33072 51708 33136 51712
rect 33072 51652 33076 51708
rect 33076 51652 33132 51708
rect 33132 51652 33136 51708
rect 33072 51648 33136 51652
rect 33152 51708 33216 51712
rect 33152 51652 33156 51708
rect 33156 51652 33212 51708
rect 33212 51652 33216 51708
rect 33152 51648 33216 51652
rect 33232 51708 33296 51712
rect 33232 51652 33236 51708
rect 33236 51652 33292 51708
rect 33292 51652 33296 51708
rect 33232 51648 33296 51652
rect 33312 51708 33376 51712
rect 33312 51652 33316 51708
rect 33316 51652 33372 51708
rect 33372 51652 33376 51708
rect 33312 51648 33376 51652
rect 3012 51164 3076 51168
rect 3012 51108 3016 51164
rect 3016 51108 3072 51164
rect 3072 51108 3076 51164
rect 3012 51104 3076 51108
rect 3092 51164 3156 51168
rect 3092 51108 3096 51164
rect 3096 51108 3152 51164
rect 3152 51108 3156 51164
rect 3092 51104 3156 51108
rect 3172 51164 3236 51168
rect 3172 51108 3176 51164
rect 3176 51108 3232 51164
rect 3232 51108 3236 51164
rect 3172 51104 3236 51108
rect 3252 51164 3316 51168
rect 3252 51108 3256 51164
rect 3256 51108 3312 51164
rect 3312 51108 3316 51164
rect 3252 51104 3316 51108
rect 33732 51164 33796 51168
rect 33732 51108 33736 51164
rect 33736 51108 33792 51164
rect 33792 51108 33796 51164
rect 33732 51104 33796 51108
rect 33812 51164 33876 51168
rect 33812 51108 33816 51164
rect 33816 51108 33872 51164
rect 33872 51108 33876 51164
rect 33812 51104 33876 51108
rect 33892 51164 33956 51168
rect 33892 51108 33896 51164
rect 33896 51108 33952 51164
rect 33952 51108 33956 51164
rect 33892 51104 33956 51108
rect 33972 51164 34036 51168
rect 33972 51108 33976 51164
rect 33976 51108 34032 51164
rect 34032 51108 34036 51164
rect 33972 51104 34036 51108
rect 2352 50620 2416 50624
rect 2352 50564 2356 50620
rect 2356 50564 2412 50620
rect 2412 50564 2416 50620
rect 2352 50560 2416 50564
rect 2432 50620 2496 50624
rect 2432 50564 2436 50620
rect 2436 50564 2492 50620
rect 2492 50564 2496 50620
rect 2432 50560 2496 50564
rect 2512 50620 2576 50624
rect 2512 50564 2516 50620
rect 2516 50564 2572 50620
rect 2572 50564 2576 50620
rect 2512 50560 2576 50564
rect 2592 50620 2656 50624
rect 2592 50564 2596 50620
rect 2596 50564 2652 50620
rect 2652 50564 2656 50620
rect 2592 50560 2656 50564
rect 33072 50620 33136 50624
rect 33072 50564 33076 50620
rect 33076 50564 33132 50620
rect 33132 50564 33136 50620
rect 33072 50560 33136 50564
rect 33152 50620 33216 50624
rect 33152 50564 33156 50620
rect 33156 50564 33212 50620
rect 33212 50564 33216 50620
rect 33152 50560 33216 50564
rect 33232 50620 33296 50624
rect 33232 50564 33236 50620
rect 33236 50564 33292 50620
rect 33292 50564 33296 50620
rect 33232 50560 33296 50564
rect 33312 50620 33376 50624
rect 33312 50564 33316 50620
rect 33316 50564 33372 50620
rect 33372 50564 33376 50620
rect 33312 50560 33376 50564
rect 3012 50076 3076 50080
rect 3012 50020 3016 50076
rect 3016 50020 3072 50076
rect 3072 50020 3076 50076
rect 3012 50016 3076 50020
rect 3092 50076 3156 50080
rect 3092 50020 3096 50076
rect 3096 50020 3152 50076
rect 3152 50020 3156 50076
rect 3092 50016 3156 50020
rect 3172 50076 3236 50080
rect 3172 50020 3176 50076
rect 3176 50020 3232 50076
rect 3232 50020 3236 50076
rect 3172 50016 3236 50020
rect 3252 50076 3316 50080
rect 3252 50020 3256 50076
rect 3256 50020 3312 50076
rect 3312 50020 3316 50076
rect 3252 50016 3316 50020
rect 33732 50076 33796 50080
rect 33732 50020 33736 50076
rect 33736 50020 33792 50076
rect 33792 50020 33796 50076
rect 33732 50016 33796 50020
rect 33812 50076 33876 50080
rect 33812 50020 33816 50076
rect 33816 50020 33872 50076
rect 33872 50020 33876 50076
rect 33812 50016 33876 50020
rect 33892 50076 33956 50080
rect 33892 50020 33896 50076
rect 33896 50020 33952 50076
rect 33952 50020 33956 50076
rect 33892 50016 33956 50020
rect 33972 50076 34036 50080
rect 33972 50020 33976 50076
rect 33976 50020 34032 50076
rect 34032 50020 34036 50076
rect 33972 50016 34036 50020
rect 2352 49532 2416 49536
rect 2352 49476 2356 49532
rect 2356 49476 2412 49532
rect 2412 49476 2416 49532
rect 2352 49472 2416 49476
rect 2432 49532 2496 49536
rect 2432 49476 2436 49532
rect 2436 49476 2492 49532
rect 2492 49476 2496 49532
rect 2432 49472 2496 49476
rect 2512 49532 2576 49536
rect 2512 49476 2516 49532
rect 2516 49476 2572 49532
rect 2572 49476 2576 49532
rect 2512 49472 2576 49476
rect 2592 49532 2656 49536
rect 2592 49476 2596 49532
rect 2596 49476 2652 49532
rect 2652 49476 2656 49532
rect 2592 49472 2656 49476
rect 33072 49532 33136 49536
rect 33072 49476 33076 49532
rect 33076 49476 33132 49532
rect 33132 49476 33136 49532
rect 33072 49472 33136 49476
rect 33152 49532 33216 49536
rect 33152 49476 33156 49532
rect 33156 49476 33212 49532
rect 33212 49476 33216 49532
rect 33152 49472 33216 49476
rect 33232 49532 33296 49536
rect 33232 49476 33236 49532
rect 33236 49476 33292 49532
rect 33292 49476 33296 49532
rect 33232 49472 33296 49476
rect 33312 49532 33376 49536
rect 33312 49476 33316 49532
rect 33316 49476 33372 49532
rect 33372 49476 33376 49532
rect 33312 49472 33376 49476
rect 3012 48988 3076 48992
rect 3012 48932 3016 48988
rect 3016 48932 3072 48988
rect 3072 48932 3076 48988
rect 3012 48928 3076 48932
rect 3092 48988 3156 48992
rect 3092 48932 3096 48988
rect 3096 48932 3152 48988
rect 3152 48932 3156 48988
rect 3092 48928 3156 48932
rect 3172 48988 3236 48992
rect 3172 48932 3176 48988
rect 3176 48932 3232 48988
rect 3232 48932 3236 48988
rect 3172 48928 3236 48932
rect 3252 48988 3316 48992
rect 3252 48932 3256 48988
rect 3256 48932 3312 48988
rect 3312 48932 3316 48988
rect 3252 48928 3316 48932
rect 33732 48988 33796 48992
rect 33732 48932 33736 48988
rect 33736 48932 33792 48988
rect 33792 48932 33796 48988
rect 33732 48928 33796 48932
rect 33812 48988 33876 48992
rect 33812 48932 33816 48988
rect 33816 48932 33872 48988
rect 33872 48932 33876 48988
rect 33812 48928 33876 48932
rect 33892 48988 33956 48992
rect 33892 48932 33896 48988
rect 33896 48932 33952 48988
rect 33952 48932 33956 48988
rect 33892 48928 33956 48932
rect 33972 48988 34036 48992
rect 33972 48932 33976 48988
rect 33976 48932 34032 48988
rect 34032 48932 34036 48988
rect 33972 48928 34036 48932
rect 2352 48444 2416 48448
rect 2352 48388 2356 48444
rect 2356 48388 2412 48444
rect 2412 48388 2416 48444
rect 2352 48384 2416 48388
rect 2432 48444 2496 48448
rect 2432 48388 2436 48444
rect 2436 48388 2492 48444
rect 2492 48388 2496 48444
rect 2432 48384 2496 48388
rect 2512 48444 2576 48448
rect 2512 48388 2516 48444
rect 2516 48388 2572 48444
rect 2572 48388 2576 48444
rect 2512 48384 2576 48388
rect 2592 48444 2656 48448
rect 2592 48388 2596 48444
rect 2596 48388 2652 48444
rect 2652 48388 2656 48444
rect 2592 48384 2656 48388
rect 33072 48444 33136 48448
rect 33072 48388 33076 48444
rect 33076 48388 33132 48444
rect 33132 48388 33136 48444
rect 33072 48384 33136 48388
rect 33152 48444 33216 48448
rect 33152 48388 33156 48444
rect 33156 48388 33212 48444
rect 33212 48388 33216 48444
rect 33152 48384 33216 48388
rect 33232 48444 33296 48448
rect 33232 48388 33236 48444
rect 33236 48388 33292 48444
rect 33292 48388 33296 48444
rect 33232 48384 33296 48388
rect 33312 48444 33376 48448
rect 33312 48388 33316 48444
rect 33316 48388 33372 48444
rect 33372 48388 33376 48444
rect 33312 48384 33376 48388
rect 3012 47900 3076 47904
rect 3012 47844 3016 47900
rect 3016 47844 3072 47900
rect 3072 47844 3076 47900
rect 3012 47840 3076 47844
rect 3092 47900 3156 47904
rect 3092 47844 3096 47900
rect 3096 47844 3152 47900
rect 3152 47844 3156 47900
rect 3092 47840 3156 47844
rect 3172 47900 3236 47904
rect 3172 47844 3176 47900
rect 3176 47844 3232 47900
rect 3232 47844 3236 47900
rect 3172 47840 3236 47844
rect 3252 47900 3316 47904
rect 3252 47844 3256 47900
rect 3256 47844 3312 47900
rect 3312 47844 3316 47900
rect 3252 47840 3316 47844
rect 33732 47900 33796 47904
rect 33732 47844 33736 47900
rect 33736 47844 33792 47900
rect 33792 47844 33796 47900
rect 33732 47840 33796 47844
rect 33812 47900 33876 47904
rect 33812 47844 33816 47900
rect 33816 47844 33872 47900
rect 33872 47844 33876 47900
rect 33812 47840 33876 47844
rect 33892 47900 33956 47904
rect 33892 47844 33896 47900
rect 33896 47844 33952 47900
rect 33952 47844 33956 47900
rect 33892 47840 33956 47844
rect 33972 47900 34036 47904
rect 33972 47844 33976 47900
rect 33976 47844 34032 47900
rect 34032 47844 34036 47900
rect 33972 47840 34036 47844
rect 2352 47356 2416 47360
rect 2352 47300 2356 47356
rect 2356 47300 2412 47356
rect 2412 47300 2416 47356
rect 2352 47296 2416 47300
rect 2432 47356 2496 47360
rect 2432 47300 2436 47356
rect 2436 47300 2492 47356
rect 2492 47300 2496 47356
rect 2432 47296 2496 47300
rect 2512 47356 2576 47360
rect 2512 47300 2516 47356
rect 2516 47300 2572 47356
rect 2572 47300 2576 47356
rect 2512 47296 2576 47300
rect 2592 47356 2656 47360
rect 2592 47300 2596 47356
rect 2596 47300 2652 47356
rect 2652 47300 2656 47356
rect 2592 47296 2656 47300
rect 33072 47356 33136 47360
rect 33072 47300 33076 47356
rect 33076 47300 33132 47356
rect 33132 47300 33136 47356
rect 33072 47296 33136 47300
rect 33152 47356 33216 47360
rect 33152 47300 33156 47356
rect 33156 47300 33212 47356
rect 33212 47300 33216 47356
rect 33152 47296 33216 47300
rect 33232 47356 33296 47360
rect 33232 47300 33236 47356
rect 33236 47300 33292 47356
rect 33292 47300 33296 47356
rect 33232 47296 33296 47300
rect 33312 47356 33376 47360
rect 33312 47300 33316 47356
rect 33316 47300 33372 47356
rect 33372 47300 33376 47356
rect 33312 47296 33376 47300
rect 3012 46812 3076 46816
rect 3012 46756 3016 46812
rect 3016 46756 3072 46812
rect 3072 46756 3076 46812
rect 3012 46752 3076 46756
rect 3092 46812 3156 46816
rect 3092 46756 3096 46812
rect 3096 46756 3152 46812
rect 3152 46756 3156 46812
rect 3092 46752 3156 46756
rect 3172 46812 3236 46816
rect 3172 46756 3176 46812
rect 3176 46756 3232 46812
rect 3232 46756 3236 46812
rect 3172 46752 3236 46756
rect 3252 46812 3316 46816
rect 3252 46756 3256 46812
rect 3256 46756 3312 46812
rect 3312 46756 3316 46812
rect 3252 46752 3316 46756
rect 33732 46812 33796 46816
rect 33732 46756 33736 46812
rect 33736 46756 33792 46812
rect 33792 46756 33796 46812
rect 33732 46752 33796 46756
rect 33812 46812 33876 46816
rect 33812 46756 33816 46812
rect 33816 46756 33872 46812
rect 33872 46756 33876 46812
rect 33812 46752 33876 46756
rect 33892 46812 33956 46816
rect 33892 46756 33896 46812
rect 33896 46756 33952 46812
rect 33952 46756 33956 46812
rect 33892 46752 33956 46756
rect 33972 46812 34036 46816
rect 33972 46756 33976 46812
rect 33976 46756 34032 46812
rect 34032 46756 34036 46812
rect 33972 46752 34036 46756
rect 2352 46268 2416 46272
rect 2352 46212 2356 46268
rect 2356 46212 2412 46268
rect 2412 46212 2416 46268
rect 2352 46208 2416 46212
rect 2432 46268 2496 46272
rect 2432 46212 2436 46268
rect 2436 46212 2492 46268
rect 2492 46212 2496 46268
rect 2432 46208 2496 46212
rect 2512 46268 2576 46272
rect 2512 46212 2516 46268
rect 2516 46212 2572 46268
rect 2572 46212 2576 46268
rect 2512 46208 2576 46212
rect 2592 46268 2656 46272
rect 2592 46212 2596 46268
rect 2596 46212 2652 46268
rect 2652 46212 2656 46268
rect 2592 46208 2656 46212
rect 33072 46268 33136 46272
rect 33072 46212 33076 46268
rect 33076 46212 33132 46268
rect 33132 46212 33136 46268
rect 33072 46208 33136 46212
rect 33152 46268 33216 46272
rect 33152 46212 33156 46268
rect 33156 46212 33212 46268
rect 33212 46212 33216 46268
rect 33152 46208 33216 46212
rect 33232 46268 33296 46272
rect 33232 46212 33236 46268
rect 33236 46212 33292 46268
rect 33292 46212 33296 46268
rect 33232 46208 33296 46212
rect 33312 46268 33376 46272
rect 33312 46212 33316 46268
rect 33316 46212 33372 46268
rect 33372 46212 33376 46268
rect 33312 46208 33376 46212
rect 3012 45724 3076 45728
rect 3012 45668 3016 45724
rect 3016 45668 3072 45724
rect 3072 45668 3076 45724
rect 3012 45664 3076 45668
rect 3092 45724 3156 45728
rect 3092 45668 3096 45724
rect 3096 45668 3152 45724
rect 3152 45668 3156 45724
rect 3092 45664 3156 45668
rect 3172 45724 3236 45728
rect 3172 45668 3176 45724
rect 3176 45668 3232 45724
rect 3232 45668 3236 45724
rect 3172 45664 3236 45668
rect 3252 45724 3316 45728
rect 3252 45668 3256 45724
rect 3256 45668 3312 45724
rect 3312 45668 3316 45724
rect 3252 45664 3316 45668
rect 33732 45724 33796 45728
rect 33732 45668 33736 45724
rect 33736 45668 33792 45724
rect 33792 45668 33796 45724
rect 33732 45664 33796 45668
rect 33812 45724 33876 45728
rect 33812 45668 33816 45724
rect 33816 45668 33872 45724
rect 33872 45668 33876 45724
rect 33812 45664 33876 45668
rect 33892 45724 33956 45728
rect 33892 45668 33896 45724
rect 33896 45668 33952 45724
rect 33952 45668 33956 45724
rect 33892 45664 33956 45668
rect 33972 45724 34036 45728
rect 33972 45668 33976 45724
rect 33976 45668 34032 45724
rect 34032 45668 34036 45724
rect 33972 45664 34036 45668
rect 2352 45180 2416 45184
rect 2352 45124 2356 45180
rect 2356 45124 2412 45180
rect 2412 45124 2416 45180
rect 2352 45120 2416 45124
rect 2432 45180 2496 45184
rect 2432 45124 2436 45180
rect 2436 45124 2492 45180
rect 2492 45124 2496 45180
rect 2432 45120 2496 45124
rect 2512 45180 2576 45184
rect 2512 45124 2516 45180
rect 2516 45124 2572 45180
rect 2572 45124 2576 45180
rect 2512 45120 2576 45124
rect 2592 45180 2656 45184
rect 2592 45124 2596 45180
rect 2596 45124 2652 45180
rect 2652 45124 2656 45180
rect 2592 45120 2656 45124
rect 33072 45180 33136 45184
rect 33072 45124 33076 45180
rect 33076 45124 33132 45180
rect 33132 45124 33136 45180
rect 33072 45120 33136 45124
rect 33152 45180 33216 45184
rect 33152 45124 33156 45180
rect 33156 45124 33212 45180
rect 33212 45124 33216 45180
rect 33152 45120 33216 45124
rect 33232 45180 33296 45184
rect 33232 45124 33236 45180
rect 33236 45124 33292 45180
rect 33292 45124 33296 45180
rect 33232 45120 33296 45124
rect 33312 45180 33376 45184
rect 33312 45124 33316 45180
rect 33316 45124 33372 45180
rect 33372 45124 33376 45180
rect 33312 45120 33376 45124
rect 3012 44636 3076 44640
rect 3012 44580 3016 44636
rect 3016 44580 3072 44636
rect 3072 44580 3076 44636
rect 3012 44576 3076 44580
rect 3092 44636 3156 44640
rect 3092 44580 3096 44636
rect 3096 44580 3152 44636
rect 3152 44580 3156 44636
rect 3092 44576 3156 44580
rect 3172 44636 3236 44640
rect 3172 44580 3176 44636
rect 3176 44580 3232 44636
rect 3232 44580 3236 44636
rect 3172 44576 3236 44580
rect 3252 44636 3316 44640
rect 3252 44580 3256 44636
rect 3256 44580 3312 44636
rect 3312 44580 3316 44636
rect 3252 44576 3316 44580
rect 33732 44636 33796 44640
rect 33732 44580 33736 44636
rect 33736 44580 33792 44636
rect 33792 44580 33796 44636
rect 33732 44576 33796 44580
rect 33812 44636 33876 44640
rect 33812 44580 33816 44636
rect 33816 44580 33872 44636
rect 33872 44580 33876 44636
rect 33812 44576 33876 44580
rect 33892 44636 33956 44640
rect 33892 44580 33896 44636
rect 33896 44580 33952 44636
rect 33952 44580 33956 44636
rect 33892 44576 33956 44580
rect 33972 44636 34036 44640
rect 33972 44580 33976 44636
rect 33976 44580 34032 44636
rect 34032 44580 34036 44636
rect 33972 44576 34036 44580
rect 2352 44092 2416 44096
rect 2352 44036 2356 44092
rect 2356 44036 2412 44092
rect 2412 44036 2416 44092
rect 2352 44032 2416 44036
rect 2432 44092 2496 44096
rect 2432 44036 2436 44092
rect 2436 44036 2492 44092
rect 2492 44036 2496 44092
rect 2432 44032 2496 44036
rect 2512 44092 2576 44096
rect 2512 44036 2516 44092
rect 2516 44036 2572 44092
rect 2572 44036 2576 44092
rect 2512 44032 2576 44036
rect 2592 44092 2656 44096
rect 2592 44036 2596 44092
rect 2596 44036 2652 44092
rect 2652 44036 2656 44092
rect 2592 44032 2656 44036
rect 33072 44092 33136 44096
rect 33072 44036 33076 44092
rect 33076 44036 33132 44092
rect 33132 44036 33136 44092
rect 33072 44032 33136 44036
rect 33152 44092 33216 44096
rect 33152 44036 33156 44092
rect 33156 44036 33212 44092
rect 33212 44036 33216 44092
rect 33152 44032 33216 44036
rect 33232 44092 33296 44096
rect 33232 44036 33236 44092
rect 33236 44036 33292 44092
rect 33292 44036 33296 44092
rect 33232 44032 33296 44036
rect 33312 44092 33376 44096
rect 33312 44036 33316 44092
rect 33316 44036 33372 44092
rect 33372 44036 33376 44092
rect 33312 44032 33376 44036
rect 3012 43548 3076 43552
rect 3012 43492 3016 43548
rect 3016 43492 3072 43548
rect 3072 43492 3076 43548
rect 3012 43488 3076 43492
rect 3092 43548 3156 43552
rect 3092 43492 3096 43548
rect 3096 43492 3152 43548
rect 3152 43492 3156 43548
rect 3092 43488 3156 43492
rect 3172 43548 3236 43552
rect 3172 43492 3176 43548
rect 3176 43492 3232 43548
rect 3232 43492 3236 43548
rect 3172 43488 3236 43492
rect 3252 43548 3316 43552
rect 3252 43492 3256 43548
rect 3256 43492 3312 43548
rect 3312 43492 3316 43548
rect 3252 43488 3316 43492
rect 33732 43548 33796 43552
rect 33732 43492 33736 43548
rect 33736 43492 33792 43548
rect 33792 43492 33796 43548
rect 33732 43488 33796 43492
rect 33812 43548 33876 43552
rect 33812 43492 33816 43548
rect 33816 43492 33872 43548
rect 33872 43492 33876 43548
rect 33812 43488 33876 43492
rect 33892 43548 33956 43552
rect 33892 43492 33896 43548
rect 33896 43492 33952 43548
rect 33952 43492 33956 43548
rect 33892 43488 33956 43492
rect 33972 43548 34036 43552
rect 33972 43492 33976 43548
rect 33976 43492 34032 43548
rect 34032 43492 34036 43548
rect 33972 43488 34036 43492
rect 2352 43004 2416 43008
rect 2352 42948 2356 43004
rect 2356 42948 2412 43004
rect 2412 42948 2416 43004
rect 2352 42944 2416 42948
rect 2432 43004 2496 43008
rect 2432 42948 2436 43004
rect 2436 42948 2492 43004
rect 2492 42948 2496 43004
rect 2432 42944 2496 42948
rect 2512 43004 2576 43008
rect 2512 42948 2516 43004
rect 2516 42948 2572 43004
rect 2572 42948 2576 43004
rect 2512 42944 2576 42948
rect 2592 43004 2656 43008
rect 2592 42948 2596 43004
rect 2596 42948 2652 43004
rect 2652 42948 2656 43004
rect 2592 42944 2656 42948
rect 33072 43004 33136 43008
rect 33072 42948 33076 43004
rect 33076 42948 33132 43004
rect 33132 42948 33136 43004
rect 33072 42944 33136 42948
rect 33152 43004 33216 43008
rect 33152 42948 33156 43004
rect 33156 42948 33212 43004
rect 33212 42948 33216 43004
rect 33152 42944 33216 42948
rect 33232 43004 33296 43008
rect 33232 42948 33236 43004
rect 33236 42948 33292 43004
rect 33292 42948 33296 43004
rect 33232 42944 33296 42948
rect 33312 43004 33376 43008
rect 33312 42948 33316 43004
rect 33316 42948 33372 43004
rect 33372 42948 33376 43004
rect 33312 42944 33376 42948
rect 3012 42460 3076 42464
rect 3012 42404 3016 42460
rect 3016 42404 3072 42460
rect 3072 42404 3076 42460
rect 3012 42400 3076 42404
rect 3092 42460 3156 42464
rect 3092 42404 3096 42460
rect 3096 42404 3152 42460
rect 3152 42404 3156 42460
rect 3092 42400 3156 42404
rect 3172 42460 3236 42464
rect 3172 42404 3176 42460
rect 3176 42404 3232 42460
rect 3232 42404 3236 42460
rect 3172 42400 3236 42404
rect 3252 42460 3316 42464
rect 3252 42404 3256 42460
rect 3256 42404 3312 42460
rect 3312 42404 3316 42460
rect 3252 42400 3316 42404
rect 33732 42460 33796 42464
rect 33732 42404 33736 42460
rect 33736 42404 33792 42460
rect 33792 42404 33796 42460
rect 33732 42400 33796 42404
rect 33812 42460 33876 42464
rect 33812 42404 33816 42460
rect 33816 42404 33872 42460
rect 33872 42404 33876 42460
rect 33812 42400 33876 42404
rect 33892 42460 33956 42464
rect 33892 42404 33896 42460
rect 33896 42404 33952 42460
rect 33952 42404 33956 42460
rect 33892 42400 33956 42404
rect 33972 42460 34036 42464
rect 33972 42404 33976 42460
rect 33976 42404 34032 42460
rect 34032 42404 34036 42460
rect 33972 42400 34036 42404
rect 2352 41916 2416 41920
rect 2352 41860 2356 41916
rect 2356 41860 2412 41916
rect 2412 41860 2416 41916
rect 2352 41856 2416 41860
rect 2432 41916 2496 41920
rect 2432 41860 2436 41916
rect 2436 41860 2492 41916
rect 2492 41860 2496 41916
rect 2432 41856 2496 41860
rect 2512 41916 2576 41920
rect 2512 41860 2516 41916
rect 2516 41860 2572 41916
rect 2572 41860 2576 41916
rect 2512 41856 2576 41860
rect 2592 41916 2656 41920
rect 2592 41860 2596 41916
rect 2596 41860 2652 41916
rect 2652 41860 2656 41916
rect 2592 41856 2656 41860
rect 33072 41916 33136 41920
rect 33072 41860 33076 41916
rect 33076 41860 33132 41916
rect 33132 41860 33136 41916
rect 33072 41856 33136 41860
rect 33152 41916 33216 41920
rect 33152 41860 33156 41916
rect 33156 41860 33212 41916
rect 33212 41860 33216 41916
rect 33152 41856 33216 41860
rect 33232 41916 33296 41920
rect 33232 41860 33236 41916
rect 33236 41860 33292 41916
rect 33292 41860 33296 41916
rect 33232 41856 33296 41860
rect 33312 41916 33376 41920
rect 33312 41860 33316 41916
rect 33316 41860 33372 41916
rect 33372 41860 33376 41916
rect 33312 41856 33376 41860
rect 3012 41372 3076 41376
rect 3012 41316 3016 41372
rect 3016 41316 3072 41372
rect 3072 41316 3076 41372
rect 3012 41312 3076 41316
rect 3092 41372 3156 41376
rect 3092 41316 3096 41372
rect 3096 41316 3152 41372
rect 3152 41316 3156 41372
rect 3092 41312 3156 41316
rect 3172 41372 3236 41376
rect 3172 41316 3176 41372
rect 3176 41316 3232 41372
rect 3232 41316 3236 41372
rect 3172 41312 3236 41316
rect 3252 41372 3316 41376
rect 3252 41316 3256 41372
rect 3256 41316 3312 41372
rect 3312 41316 3316 41372
rect 3252 41312 3316 41316
rect 33732 41372 33796 41376
rect 33732 41316 33736 41372
rect 33736 41316 33792 41372
rect 33792 41316 33796 41372
rect 33732 41312 33796 41316
rect 33812 41372 33876 41376
rect 33812 41316 33816 41372
rect 33816 41316 33872 41372
rect 33872 41316 33876 41372
rect 33812 41312 33876 41316
rect 33892 41372 33956 41376
rect 33892 41316 33896 41372
rect 33896 41316 33952 41372
rect 33952 41316 33956 41372
rect 33892 41312 33956 41316
rect 33972 41372 34036 41376
rect 33972 41316 33976 41372
rect 33976 41316 34032 41372
rect 34032 41316 34036 41372
rect 33972 41312 34036 41316
rect 2352 40828 2416 40832
rect 2352 40772 2356 40828
rect 2356 40772 2412 40828
rect 2412 40772 2416 40828
rect 2352 40768 2416 40772
rect 2432 40828 2496 40832
rect 2432 40772 2436 40828
rect 2436 40772 2492 40828
rect 2492 40772 2496 40828
rect 2432 40768 2496 40772
rect 2512 40828 2576 40832
rect 2512 40772 2516 40828
rect 2516 40772 2572 40828
rect 2572 40772 2576 40828
rect 2512 40768 2576 40772
rect 2592 40828 2656 40832
rect 2592 40772 2596 40828
rect 2596 40772 2652 40828
rect 2652 40772 2656 40828
rect 2592 40768 2656 40772
rect 33072 40828 33136 40832
rect 33072 40772 33076 40828
rect 33076 40772 33132 40828
rect 33132 40772 33136 40828
rect 33072 40768 33136 40772
rect 33152 40828 33216 40832
rect 33152 40772 33156 40828
rect 33156 40772 33212 40828
rect 33212 40772 33216 40828
rect 33152 40768 33216 40772
rect 33232 40828 33296 40832
rect 33232 40772 33236 40828
rect 33236 40772 33292 40828
rect 33292 40772 33296 40828
rect 33232 40768 33296 40772
rect 33312 40828 33376 40832
rect 33312 40772 33316 40828
rect 33316 40772 33372 40828
rect 33372 40772 33376 40828
rect 33312 40768 33376 40772
rect 3012 40284 3076 40288
rect 3012 40228 3016 40284
rect 3016 40228 3072 40284
rect 3072 40228 3076 40284
rect 3012 40224 3076 40228
rect 3092 40284 3156 40288
rect 3092 40228 3096 40284
rect 3096 40228 3152 40284
rect 3152 40228 3156 40284
rect 3092 40224 3156 40228
rect 3172 40284 3236 40288
rect 3172 40228 3176 40284
rect 3176 40228 3232 40284
rect 3232 40228 3236 40284
rect 3172 40224 3236 40228
rect 3252 40284 3316 40288
rect 3252 40228 3256 40284
rect 3256 40228 3312 40284
rect 3312 40228 3316 40284
rect 3252 40224 3316 40228
rect 33732 40284 33796 40288
rect 33732 40228 33736 40284
rect 33736 40228 33792 40284
rect 33792 40228 33796 40284
rect 33732 40224 33796 40228
rect 33812 40284 33876 40288
rect 33812 40228 33816 40284
rect 33816 40228 33872 40284
rect 33872 40228 33876 40284
rect 33812 40224 33876 40228
rect 33892 40284 33956 40288
rect 33892 40228 33896 40284
rect 33896 40228 33952 40284
rect 33952 40228 33956 40284
rect 33892 40224 33956 40228
rect 33972 40284 34036 40288
rect 33972 40228 33976 40284
rect 33976 40228 34032 40284
rect 34032 40228 34036 40284
rect 33972 40224 34036 40228
rect 2352 39740 2416 39744
rect 2352 39684 2356 39740
rect 2356 39684 2412 39740
rect 2412 39684 2416 39740
rect 2352 39680 2416 39684
rect 2432 39740 2496 39744
rect 2432 39684 2436 39740
rect 2436 39684 2492 39740
rect 2492 39684 2496 39740
rect 2432 39680 2496 39684
rect 2512 39740 2576 39744
rect 2512 39684 2516 39740
rect 2516 39684 2572 39740
rect 2572 39684 2576 39740
rect 2512 39680 2576 39684
rect 2592 39740 2656 39744
rect 2592 39684 2596 39740
rect 2596 39684 2652 39740
rect 2652 39684 2656 39740
rect 2592 39680 2656 39684
rect 33072 39740 33136 39744
rect 33072 39684 33076 39740
rect 33076 39684 33132 39740
rect 33132 39684 33136 39740
rect 33072 39680 33136 39684
rect 33152 39740 33216 39744
rect 33152 39684 33156 39740
rect 33156 39684 33212 39740
rect 33212 39684 33216 39740
rect 33152 39680 33216 39684
rect 33232 39740 33296 39744
rect 33232 39684 33236 39740
rect 33236 39684 33292 39740
rect 33292 39684 33296 39740
rect 33232 39680 33296 39684
rect 33312 39740 33376 39744
rect 33312 39684 33316 39740
rect 33316 39684 33372 39740
rect 33372 39684 33376 39740
rect 33312 39680 33376 39684
rect 3012 39196 3076 39200
rect 3012 39140 3016 39196
rect 3016 39140 3072 39196
rect 3072 39140 3076 39196
rect 3012 39136 3076 39140
rect 3092 39196 3156 39200
rect 3092 39140 3096 39196
rect 3096 39140 3152 39196
rect 3152 39140 3156 39196
rect 3092 39136 3156 39140
rect 3172 39196 3236 39200
rect 3172 39140 3176 39196
rect 3176 39140 3232 39196
rect 3232 39140 3236 39196
rect 3172 39136 3236 39140
rect 3252 39196 3316 39200
rect 3252 39140 3256 39196
rect 3256 39140 3312 39196
rect 3312 39140 3316 39196
rect 3252 39136 3316 39140
rect 33732 39196 33796 39200
rect 33732 39140 33736 39196
rect 33736 39140 33792 39196
rect 33792 39140 33796 39196
rect 33732 39136 33796 39140
rect 33812 39196 33876 39200
rect 33812 39140 33816 39196
rect 33816 39140 33872 39196
rect 33872 39140 33876 39196
rect 33812 39136 33876 39140
rect 33892 39196 33956 39200
rect 33892 39140 33896 39196
rect 33896 39140 33952 39196
rect 33952 39140 33956 39196
rect 33892 39136 33956 39140
rect 33972 39196 34036 39200
rect 33972 39140 33976 39196
rect 33976 39140 34032 39196
rect 34032 39140 34036 39196
rect 33972 39136 34036 39140
rect 2352 38652 2416 38656
rect 2352 38596 2356 38652
rect 2356 38596 2412 38652
rect 2412 38596 2416 38652
rect 2352 38592 2416 38596
rect 2432 38652 2496 38656
rect 2432 38596 2436 38652
rect 2436 38596 2492 38652
rect 2492 38596 2496 38652
rect 2432 38592 2496 38596
rect 2512 38652 2576 38656
rect 2512 38596 2516 38652
rect 2516 38596 2572 38652
rect 2572 38596 2576 38652
rect 2512 38592 2576 38596
rect 2592 38652 2656 38656
rect 2592 38596 2596 38652
rect 2596 38596 2652 38652
rect 2652 38596 2656 38652
rect 2592 38592 2656 38596
rect 33072 38652 33136 38656
rect 33072 38596 33076 38652
rect 33076 38596 33132 38652
rect 33132 38596 33136 38652
rect 33072 38592 33136 38596
rect 33152 38652 33216 38656
rect 33152 38596 33156 38652
rect 33156 38596 33212 38652
rect 33212 38596 33216 38652
rect 33152 38592 33216 38596
rect 33232 38652 33296 38656
rect 33232 38596 33236 38652
rect 33236 38596 33292 38652
rect 33292 38596 33296 38652
rect 33232 38592 33296 38596
rect 33312 38652 33376 38656
rect 33312 38596 33316 38652
rect 33316 38596 33372 38652
rect 33372 38596 33376 38652
rect 33312 38592 33376 38596
rect 3012 38108 3076 38112
rect 3012 38052 3016 38108
rect 3016 38052 3072 38108
rect 3072 38052 3076 38108
rect 3012 38048 3076 38052
rect 3092 38108 3156 38112
rect 3092 38052 3096 38108
rect 3096 38052 3152 38108
rect 3152 38052 3156 38108
rect 3092 38048 3156 38052
rect 3172 38108 3236 38112
rect 3172 38052 3176 38108
rect 3176 38052 3232 38108
rect 3232 38052 3236 38108
rect 3172 38048 3236 38052
rect 3252 38108 3316 38112
rect 3252 38052 3256 38108
rect 3256 38052 3312 38108
rect 3312 38052 3316 38108
rect 3252 38048 3316 38052
rect 33732 38108 33796 38112
rect 33732 38052 33736 38108
rect 33736 38052 33792 38108
rect 33792 38052 33796 38108
rect 33732 38048 33796 38052
rect 33812 38108 33876 38112
rect 33812 38052 33816 38108
rect 33816 38052 33872 38108
rect 33872 38052 33876 38108
rect 33812 38048 33876 38052
rect 33892 38108 33956 38112
rect 33892 38052 33896 38108
rect 33896 38052 33952 38108
rect 33952 38052 33956 38108
rect 33892 38048 33956 38052
rect 33972 38108 34036 38112
rect 33972 38052 33976 38108
rect 33976 38052 34032 38108
rect 34032 38052 34036 38108
rect 33972 38048 34036 38052
rect 2352 37564 2416 37568
rect 2352 37508 2356 37564
rect 2356 37508 2412 37564
rect 2412 37508 2416 37564
rect 2352 37504 2416 37508
rect 2432 37564 2496 37568
rect 2432 37508 2436 37564
rect 2436 37508 2492 37564
rect 2492 37508 2496 37564
rect 2432 37504 2496 37508
rect 2512 37564 2576 37568
rect 2512 37508 2516 37564
rect 2516 37508 2572 37564
rect 2572 37508 2576 37564
rect 2512 37504 2576 37508
rect 2592 37564 2656 37568
rect 2592 37508 2596 37564
rect 2596 37508 2652 37564
rect 2652 37508 2656 37564
rect 2592 37504 2656 37508
rect 33072 37564 33136 37568
rect 33072 37508 33076 37564
rect 33076 37508 33132 37564
rect 33132 37508 33136 37564
rect 33072 37504 33136 37508
rect 33152 37564 33216 37568
rect 33152 37508 33156 37564
rect 33156 37508 33212 37564
rect 33212 37508 33216 37564
rect 33152 37504 33216 37508
rect 33232 37564 33296 37568
rect 33232 37508 33236 37564
rect 33236 37508 33292 37564
rect 33292 37508 33296 37564
rect 33232 37504 33296 37508
rect 33312 37564 33376 37568
rect 33312 37508 33316 37564
rect 33316 37508 33372 37564
rect 33372 37508 33376 37564
rect 33312 37504 33376 37508
rect 3012 37020 3076 37024
rect 3012 36964 3016 37020
rect 3016 36964 3072 37020
rect 3072 36964 3076 37020
rect 3012 36960 3076 36964
rect 3092 37020 3156 37024
rect 3092 36964 3096 37020
rect 3096 36964 3152 37020
rect 3152 36964 3156 37020
rect 3092 36960 3156 36964
rect 3172 37020 3236 37024
rect 3172 36964 3176 37020
rect 3176 36964 3232 37020
rect 3232 36964 3236 37020
rect 3172 36960 3236 36964
rect 3252 37020 3316 37024
rect 3252 36964 3256 37020
rect 3256 36964 3312 37020
rect 3312 36964 3316 37020
rect 3252 36960 3316 36964
rect 33732 37020 33796 37024
rect 33732 36964 33736 37020
rect 33736 36964 33792 37020
rect 33792 36964 33796 37020
rect 33732 36960 33796 36964
rect 33812 37020 33876 37024
rect 33812 36964 33816 37020
rect 33816 36964 33872 37020
rect 33872 36964 33876 37020
rect 33812 36960 33876 36964
rect 33892 37020 33956 37024
rect 33892 36964 33896 37020
rect 33896 36964 33952 37020
rect 33952 36964 33956 37020
rect 33892 36960 33956 36964
rect 33972 37020 34036 37024
rect 33972 36964 33976 37020
rect 33976 36964 34032 37020
rect 34032 36964 34036 37020
rect 33972 36960 34036 36964
rect 2352 36476 2416 36480
rect 2352 36420 2356 36476
rect 2356 36420 2412 36476
rect 2412 36420 2416 36476
rect 2352 36416 2416 36420
rect 2432 36476 2496 36480
rect 2432 36420 2436 36476
rect 2436 36420 2492 36476
rect 2492 36420 2496 36476
rect 2432 36416 2496 36420
rect 2512 36476 2576 36480
rect 2512 36420 2516 36476
rect 2516 36420 2572 36476
rect 2572 36420 2576 36476
rect 2512 36416 2576 36420
rect 2592 36476 2656 36480
rect 2592 36420 2596 36476
rect 2596 36420 2652 36476
rect 2652 36420 2656 36476
rect 2592 36416 2656 36420
rect 33072 36476 33136 36480
rect 33072 36420 33076 36476
rect 33076 36420 33132 36476
rect 33132 36420 33136 36476
rect 33072 36416 33136 36420
rect 33152 36476 33216 36480
rect 33152 36420 33156 36476
rect 33156 36420 33212 36476
rect 33212 36420 33216 36476
rect 33152 36416 33216 36420
rect 33232 36476 33296 36480
rect 33232 36420 33236 36476
rect 33236 36420 33292 36476
rect 33292 36420 33296 36476
rect 33232 36416 33296 36420
rect 33312 36476 33376 36480
rect 33312 36420 33316 36476
rect 33316 36420 33372 36476
rect 33372 36420 33376 36476
rect 33312 36416 33376 36420
rect 3012 35932 3076 35936
rect 3012 35876 3016 35932
rect 3016 35876 3072 35932
rect 3072 35876 3076 35932
rect 3012 35872 3076 35876
rect 3092 35932 3156 35936
rect 3092 35876 3096 35932
rect 3096 35876 3152 35932
rect 3152 35876 3156 35932
rect 3092 35872 3156 35876
rect 3172 35932 3236 35936
rect 3172 35876 3176 35932
rect 3176 35876 3232 35932
rect 3232 35876 3236 35932
rect 3172 35872 3236 35876
rect 3252 35932 3316 35936
rect 3252 35876 3256 35932
rect 3256 35876 3312 35932
rect 3312 35876 3316 35932
rect 3252 35872 3316 35876
rect 33732 35932 33796 35936
rect 33732 35876 33736 35932
rect 33736 35876 33792 35932
rect 33792 35876 33796 35932
rect 33732 35872 33796 35876
rect 33812 35932 33876 35936
rect 33812 35876 33816 35932
rect 33816 35876 33872 35932
rect 33872 35876 33876 35932
rect 33812 35872 33876 35876
rect 33892 35932 33956 35936
rect 33892 35876 33896 35932
rect 33896 35876 33952 35932
rect 33952 35876 33956 35932
rect 33892 35872 33956 35876
rect 33972 35932 34036 35936
rect 33972 35876 33976 35932
rect 33976 35876 34032 35932
rect 34032 35876 34036 35932
rect 33972 35872 34036 35876
rect 2352 35388 2416 35392
rect 2352 35332 2356 35388
rect 2356 35332 2412 35388
rect 2412 35332 2416 35388
rect 2352 35328 2416 35332
rect 2432 35388 2496 35392
rect 2432 35332 2436 35388
rect 2436 35332 2492 35388
rect 2492 35332 2496 35388
rect 2432 35328 2496 35332
rect 2512 35388 2576 35392
rect 2512 35332 2516 35388
rect 2516 35332 2572 35388
rect 2572 35332 2576 35388
rect 2512 35328 2576 35332
rect 2592 35388 2656 35392
rect 2592 35332 2596 35388
rect 2596 35332 2652 35388
rect 2652 35332 2656 35388
rect 2592 35328 2656 35332
rect 33072 35388 33136 35392
rect 33072 35332 33076 35388
rect 33076 35332 33132 35388
rect 33132 35332 33136 35388
rect 33072 35328 33136 35332
rect 33152 35388 33216 35392
rect 33152 35332 33156 35388
rect 33156 35332 33212 35388
rect 33212 35332 33216 35388
rect 33152 35328 33216 35332
rect 33232 35388 33296 35392
rect 33232 35332 33236 35388
rect 33236 35332 33292 35388
rect 33292 35332 33296 35388
rect 33232 35328 33296 35332
rect 33312 35388 33376 35392
rect 33312 35332 33316 35388
rect 33316 35332 33372 35388
rect 33372 35332 33376 35388
rect 33312 35328 33376 35332
rect 3012 34844 3076 34848
rect 3012 34788 3016 34844
rect 3016 34788 3072 34844
rect 3072 34788 3076 34844
rect 3012 34784 3076 34788
rect 3092 34844 3156 34848
rect 3092 34788 3096 34844
rect 3096 34788 3152 34844
rect 3152 34788 3156 34844
rect 3092 34784 3156 34788
rect 3172 34844 3236 34848
rect 3172 34788 3176 34844
rect 3176 34788 3232 34844
rect 3232 34788 3236 34844
rect 3172 34784 3236 34788
rect 3252 34844 3316 34848
rect 3252 34788 3256 34844
rect 3256 34788 3312 34844
rect 3312 34788 3316 34844
rect 3252 34784 3316 34788
rect 33732 34844 33796 34848
rect 33732 34788 33736 34844
rect 33736 34788 33792 34844
rect 33792 34788 33796 34844
rect 33732 34784 33796 34788
rect 33812 34844 33876 34848
rect 33812 34788 33816 34844
rect 33816 34788 33872 34844
rect 33872 34788 33876 34844
rect 33812 34784 33876 34788
rect 33892 34844 33956 34848
rect 33892 34788 33896 34844
rect 33896 34788 33952 34844
rect 33952 34788 33956 34844
rect 33892 34784 33956 34788
rect 33972 34844 34036 34848
rect 33972 34788 33976 34844
rect 33976 34788 34032 34844
rect 34032 34788 34036 34844
rect 33972 34784 34036 34788
rect 2352 34300 2416 34304
rect 2352 34244 2356 34300
rect 2356 34244 2412 34300
rect 2412 34244 2416 34300
rect 2352 34240 2416 34244
rect 2432 34300 2496 34304
rect 2432 34244 2436 34300
rect 2436 34244 2492 34300
rect 2492 34244 2496 34300
rect 2432 34240 2496 34244
rect 2512 34300 2576 34304
rect 2512 34244 2516 34300
rect 2516 34244 2572 34300
rect 2572 34244 2576 34300
rect 2512 34240 2576 34244
rect 2592 34300 2656 34304
rect 2592 34244 2596 34300
rect 2596 34244 2652 34300
rect 2652 34244 2656 34300
rect 2592 34240 2656 34244
rect 33072 34300 33136 34304
rect 33072 34244 33076 34300
rect 33076 34244 33132 34300
rect 33132 34244 33136 34300
rect 33072 34240 33136 34244
rect 33152 34300 33216 34304
rect 33152 34244 33156 34300
rect 33156 34244 33212 34300
rect 33212 34244 33216 34300
rect 33152 34240 33216 34244
rect 33232 34300 33296 34304
rect 33232 34244 33236 34300
rect 33236 34244 33292 34300
rect 33292 34244 33296 34300
rect 33232 34240 33296 34244
rect 33312 34300 33376 34304
rect 33312 34244 33316 34300
rect 33316 34244 33372 34300
rect 33372 34244 33376 34300
rect 33312 34240 33376 34244
rect 3012 33756 3076 33760
rect 3012 33700 3016 33756
rect 3016 33700 3072 33756
rect 3072 33700 3076 33756
rect 3012 33696 3076 33700
rect 3092 33756 3156 33760
rect 3092 33700 3096 33756
rect 3096 33700 3152 33756
rect 3152 33700 3156 33756
rect 3092 33696 3156 33700
rect 3172 33756 3236 33760
rect 3172 33700 3176 33756
rect 3176 33700 3232 33756
rect 3232 33700 3236 33756
rect 3172 33696 3236 33700
rect 3252 33756 3316 33760
rect 3252 33700 3256 33756
rect 3256 33700 3312 33756
rect 3312 33700 3316 33756
rect 3252 33696 3316 33700
rect 33732 33756 33796 33760
rect 33732 33700 33736 33756
rect 33736 33700 33792 33756
rect 33792 33700 33796 33756
rect 33732 33696 33796 33700
rect 33812 33756 33876 33760
rect 33812 33700 33816 33756
rect 33816 33700 33872 33756
rect 33872 33700 33876 33756
rect 33812 33696 33876 33700
rect 33892 33756 33956 33760
rect 33892 33700 33896 33756
rect 33896 33700 33952 33756
rect 33952 33700 33956 33756
rect 33892 33696 33956 33700
rect 33972 33756 34036 33760
rect 33972 33700 33976 33756
rect 33976 33700 34032 33756
rect 34032 33700 34036 33756
rect 33972 33696 34036 33700
rect 2352 33212 2416 33216
rect 2352 33156 2356 33212
rect 2356 33156 2412 33212
rect 2412 33156 2416 33212
rect 2352 33152 2416 33156
rect 2432 33212 2496 33216
rect 2432 33156 2436 33212
rect 2436 33156 2492 33212
rect 2492 33156 2496 33212
rect 2432 33152 2496 33156
rect 2512 33212 2576 33216
rect 2512 33156 2516 33212
rect 2516 33156 2572 33212
rect 2572 33156 2576 33212
rect 2512 33152 2576 33156
rect 2592 33212 2656 33216
rect 2592 33156 2596 33212
rect 2596 33156 2652 33212
rect 2652 33156 2656 33212
rect 2592 33152 2656 33156
rect 33072 33212 33136 33216
rect 33072 33156 33076 33212
rect 33076 33156 33132 33212
rect 33132 33156 33136 33212
rect 33072 33152 33136 33156
rect 33152 33212 33216 33216
rect 33152 33156 33156 33212
rect 33156 33156 33212 33212
rect 33212 33156 33216 33212
rect 33152 33152 33216 33156
rect 33232 33212 33296 33216
rect 33232 33156 33236 33212
rect 33236 33156 33292 33212
rect 33292 33156 33296 33212
rect 33232 33152 33296 33156
rect 33312 33212 33376 33216
rect 33312 33156 33316 33212
rect 33316 33156 33372 33212
rect 33372 33156 33376 33212
rect 33312 33152 33376 33156
rect 3012 32668 3076 32672
rect 3012 32612 3016 32668
rect 3016 32612 3072 32668
rect 3072 32612 3076 32668
rect 3012 32608 3076 32612
rect 3092 32668 3156 32672
rect 3092 32612 3096 32668
rect 3096 32612 3152 32668
rect 3152 32612 3156 32668
rect 3092 32608 3156 32612
rect 3172 32668 3236 32672
rect 3172 32612 3176 32668
rect 3176 32612 3232 32668
rect 3232 32612 3236 32668
rect 3172 32608 3236 32612
rect 3252 32668 3316 32672
rect 3252 32612 3256 32668
rect 3256 32612 3312 32668
rect 3312 32612 3316 32668
rect 3252 32608 3316 32612
rect 33732 32668 33796 32672
rect 33732 32612 33736 32668
rect 33736 32612 33792 32668
rect 33792 32612 33796 32668
rect 33732 32608 33796 32612
rect 33812 32668 33876 32672
rect 33812 32612 33816 32668
rect 33816 32612 33872 32668
rect 33872 32612 33876 32668
rect 33812 32608 33876 32612
rect 33892 32668 33956 32672
rect 33892 32612 33896 32668
rect 33896 32612 33952 32668
rect 33952 32612 33956 32668
rect 33892 32608 33956 32612
rect 33972 32668 34036 32672
rect 33972 32612 33976 32668
rect 33976 32612 34032 32668
rect 34032 32612 34036 32668
rect 33972 32608 34036 32612
rect 2352 32124 2416 32128
rect 2352 32068 2356 32124
rect 2356 32068 2412 32124
rect 2412 32068 2416 32124
rect 2352 32064 2416 32068
rect 2432 32124 2496 32128
rect 2432 32068 2436 32124
rect 2436 32068 2492 32124
rect 2492 32068 2496 32124
rect 2432 32064 2496 32068
rect 2512 32124 2576 32128
rect 2512 32068 2516 32124
rect 2516 32068 2572 32124
rect 2572 32068 2576 32124
rect 2512 32064 2576 32068
rect 2592 32124 2656 32128
rect 2592 32068 2596 32124
rect 2596 32068 2652 32124
rect 2652 32068 2656 32124
rect 2592 32064 2656 32068
rect 33072 32124 33136 32128
rect 33072 32068 33076 32124
rect 33076 32068 33132 32124
rect 33132 32068 33136 32124
rect 33072 32064 33136 32068
rect 33152 32124 33216 32128
rect 33152 32068 33156 32124
rect 33156 32068 33212 32124
rect 33212 32068 33216 32124
rect 33152 32064 33216 32068
rect 33232 32124 33296 32128
rect 33232 32068 33236 32124
rect 33236 32068 33292 32124
rect 33292 32068 33296 32124
rect 33232 32064 33296 32068
rect 33312 32124 33376 32128
rect 33312 32068 33316 32124
rect 33316 32068 33372 32124
rect 33372 32068 33376 32124
rect 33312 32064 33376 32068
rect 3012 31580 3076 31584
rect 3012 31524 3016 31580
rect 3016 31524 3072 31580
rect 3072 31524 3076 31580
rect 3012 31520 3076 31524
rect 3092 31580 3156 31584
rect 3092 31524 3096 31580
rect 3096 31524 3152 31580
rect 3152 31524 3156 31580
rect 3092 31520 3156 31524
rect 3172 31580 3236 31584
rect 3172 31524 3176 31580
rect 3176 31524 3232 31580
rect 3232 31524 3236 31580
rect 3172 31520 3236 31524
rect 3252 31580 3316 31584
rect 3252 31524 3256 31580
rect 3256 31524 3312 31580
rect 3312 31524 3316 31580
rect 3252 31520 3316 31524
rect 33732 31580 33796 31584
rect 33732 31524 33736 31580
rect 33736 31524 33792 31580
rect 33792 31524 33796 31580
rect 33732 31520 33796 31524
rect 33812 31580 33876 31584
rect 33812 31524 33816 31580
rect 33816 31524 33872 31580
rect 33872 31524 33876 31580
rect 33812 31520 33876 31524
rect 33892 31580 33956 31584
rect 33892 31524 33896 31580
rect 33896 31524 33952 31580
rect 33952 31524 33956 31580
rect 33892 31520 33956 31524
rect 33972 31580 34036 31584
rect 33972 31524 33976 31580
rect 33976 31524 34032 31580
rect 34032 31524 34036 31580
rect 33972 31520 34036 31524
rect 2352 31036 2416 31040
rect 2352 30980 2356 31036
rect 2356 30980 2412 31036
rect 2412 30980 2416 31036
rect 2352 30976 2416 30980
rect 2432 31036 2496 31040
rect 2432 30980 2436 31036
rect 2436 30980 2492 31036
rect 2492 30980 2496 31036
rect 2432 30976 2496 30980
rect 2512 31036 2576 31040
rect 2512 30980 2516 31036
rect 2516 30980 2572 31036
rect 2572 30980 2576 31036
rect 2512 30976 2576 30980
rect 2592 31036 2656 31040
rect 2592 30980 2596 31036
rect 2596 30980 2652 31036
rect 2652 30980 2656 31036
rect 2592 30976 2656 30980
rect 33072 31036 33136 31040
rect 33072 30980 33076 31036
rect 33076 30980 33132 31036
rect 33132 30980 33136 31036
rect 33072 30976 33136 30980
rect 33152 31036 33216 31040
rect 33152 30980 33156 31036
rect 33156 30980 33212 31036
rect 33212 30980 33216 31036
rect 33152 30976 33216 30980
rect 33232 31036 33296 31040
rect 33232 30980 33236 31036
rect 33236 30980 33292 31036
rect 33292 30980 33296 31036
rect 33232 30976 33296 30980
rect 33312 31036 33376 31040
rect 33312 30980 33316 31036
rect 33316 30980 33372 31036
rect 33372 30980 33376 31036
rect 33312 30976 33376 30980
rect 3012 30492 3076 30496
rect 3012 30436 3016 30492
rect 3016 30436 3072 30492
rect 3072 30436 3076 30492
rect 3012 30432 3076 30436
rect 3092 30492 3156 30496
rect 3092 30436 3096 30492
rect 3096 30436 3152 30492
rect 3152 30436 3156 30492
rect 3092 30432 3156 30436
rect 3172 30492 3236 30496
rect 3172 30436 3176 30492
rect 3176 30436 3232 30492
rect 3232 30436 3236 30492
rect 3172 30432 3236 30436
rect 3252 30492 3316 30496
rect 3252 30436 3256 30492
rect 3256 30436 3312 30492
rect 3312 30436 3316 30492
rect 3252 30432 3316 30436
rect 33732 30492 33796 30496
rect 33732 30436 33736 30492
rect 33736 30436 33792 30492
rect 33792 30436 33796 30492
rect 33732 30432 33796 30436
rect 33812 30492 33876 30496
rect 33812 30436 33816 30492
rect 33816 30436 33872 30492
rect 33872 30436 33876 30492
rect 33812 30432 33876 30436
rect 33892 30492 33956 30496
rect 33892 30436 33896 30492
rect 33896 30436 33952 30492
rect 33952 30436 33956 30492
rect 33892 30432 33956 30436
rect 33972 30492 34036 30496
rect 33972 30436 33976 30492
rect 33976 30436 34032 30492
rect 34032 30436 34036 30492
rect 33972 30432 34036 30436
rect 2352 29948 2416 29952
rect 2352 29892 2356 29948
rect 2356 29892 2412 29948
rect 2412 29892 2416 29948
rect 2352 29888 2416 29892
rect 2432 29948 2496 29952
rect 2432 29892 2436 29948
rect 2436 29892 2492 29948
rect 2492 29892 2496 29948
rect 2432 29888 2496 29892
rect 2512 29948 2576 29952
rect 2512 29892 2516 29948
rect 2516 29892 2572 29948
rect 2572 29892 2576 29948
rect 2512 29888 2576 29892
rect 2592 29948 2656 29952
rect 2592 29892 2596 29948
rect 2596 29892 2652 29948
rect 2652 29892 2656 29948
rect 2592 29888 2656 29892
rect 33072 29948 33136 29952
rect 33072 29892 33076 29948
rect 33076 29892 33132 29948
rect 33132 29892 33136 29948
rect 33072 29888 33136 29892
rect 33152 29948 33216 29952
rect 33152 29892 33156 29948
rect 33156 29892 33212 29948
rect 33212 29892 33216 29948
rect 33152 29888 33216 29892
rect 33232 29948 33296 29952
rect 33232 29892 33236 29948
rect 33236 29892 33292 29948
rect 33292 29892 33296 29948
rect 33232 29888 33296 29892
rect 33312 29948 33376 29952
rect 33312 29892 33316 29948
rect 33316 29892 33372 29948
rect 33372 29892 33376 29948
rect 33312 29888 33376 29892
rect 3012 29404 3076 29408
rect 3012 29348 3016 29404
rect 3016 29348 3072 29404
rect 3072 29348 3076 29404
rect 3012 29344 3076 29348
rect 3092 29404 3156 29408
rect 3092 29348 3096 29404
rect 3096 29348 3152 29404
rect 3152 29348 3156 29404
rect 3092 29344 3156 29348
rect 3172 29404 3236 29408
rect 3172 29348 3176 29404
rect 3176 29348 3232 29404
rect 3232 29348 3236 29404
rect 3172 29344 3236 29348
rect 3252 29404 3316 29408
rect 3252 29348 3256 29404
rect 3256 29348 3312 29404
rect 3312 29348 3316 29404
rect 3252 29344 3316 29348
rect 33732 29404 33796 29408
rect 33732 29348 33736 29404
rect 33736 29348 33792 29404
rect 33792 29348 33796 29404
rect 33732 29344 33796 29348
rect 33812 29404 33876 29408
rect 33812 29348 33816 29404
rect 33816 29348 33872 29404
rect 33872 29348 33876 29404
rect 33812 29344 33876 29348
rect 33892 29404 33956 29408
rect 33892 29348 33896 29404
rect 33896 29348 33952 29404
rect 33952 29348 33956 29404
rect 33892 29344 33956 29348
rect 33972 29404 34036 29408
rect 33972 29348 33976 29404
rect 33976 29348 34032 29404
rect 34032 29348 34036 29404
rect 33972 29344 34036 29348
rect 2352 28860 2416 28864
rect 2352 28804 2356 28860
rect 2356 28804 2412 28860
rect 2412 28804 2416 28860
rect 2352 28800 2416 28804
rect 2432 28860 2496 28864
rect 2432 28804 2436 28860
rect 2436 28804 2492 28860
rect 2492 28804 2496 28860
rect 2432 28800 2496 28804
rect 2512 28860 2576 28864
rect 2512 28804 2516 28860
rect 2516 28804 2572 28860
rect 2572 28804 2576 28860
rect 2512 28800 2576 28804
rect 2592 28860 2656 28864
rect 2592 28804 2596 28860
rect 2596 28804 2652 28860
rect 2652 28804 2656 28860
rect 2592 28800 2656 28804
rect 33072 28860 33136 28864
rect 33072 28804 33076 28860
rect 33076 28804 33132 28860
rect 33132 28804 33136 28860
rect 33072 28800 33136 28804
rect 33152 28860 33216 28864
rect 33152 28804 33156 28860
rect 33156 28804 33212 28860
rect 33212 28804 33216 28860
rect 33152 28800 33216 28804
rect 33232 28860 33296 28864
rect 33232 28804 33236 28860
rect 33236 28804 33292 28860
rect 33292 28804 33296 28860
rect 33232 28800 33296 28804
rect 33312 28860 33376 28864
rect 33312 28804 33316 28860
rect 33316 28804 33372 28860
rect 33372 28804 33376 28860
rect 33312 28800 33376 28804
rect 3012 28316 3076 28320
rect 3012 28260 3016 28316
rect 3016 28260 3072 28316
rect 3072 28260 3076 28316
rect 3012 28256 3076 28260
rect 3092 28316 3156 28320
rect 3092 28260 3096 28316
rect 3096 28260 3152 28316
rect 3152 28260 3156 28316
rect 3092 28256 3156 28260
rect 3172 28316 3236 28320
rect 3172 28260 3176 28316
rect 3176 28260 3232 28316
rect 3232 28260 3236 28316
rect 3172 28256 3236 28260
rect 3252 28316 3316 28320
rect 3252 28260 3256 28316
rect 3256 28260 3312 28316
rect 3312 28260 3316 28316
rect 3252 28256 3316 28260
rect 33732 28316 33796 28320
rect 33732 28260 33736 28316
rect 33736 28260 33792 28316
rect 33792 28260 33796 28316
rect 33732 28256 33796 28260
rect 33812 28316 33876 28320
rect 33812 28260 33816 28316
rect 33816 28260 33872 28316
rect 33872 28260 33876 28316
rect 33812 28256 33876 28260
rect 33892 28316 33956 28320
rect 33892 28260 33896 28316
rect 33896 28260 33952 28316
rect 33952 28260 33956 28316
rect 33892 28256 33956 28260
rect 33972 28316 34036 28320
rect 33972 28260 33976 28316
rect 33976 28260 34032 28316
rect 34032 28260 34036 28316
rect 33972 28256 34036 28260
rect 2352 27772 2416 27776
rect 2352 27716 2356 27772
rect 2356 27716 2412 27772
rect 2412 27716 2416 27772
rect 2352 27712 2416 27716
rect 2432 27772 2496 27776
rect 2432 27716 2436 27772
rect 2436 27716 2492 27772
rect 2492 27716 2496 27772
rect 2432 27712 2496 27716
rect 2512 27772 2576 27776
rect 2512 27716 2516 27772
rect 2516 27716 2572 27772
rect 2572 27716 2576 27772
rect 2512 27712 2576 27716
rect 2592 27772 2656 27776
rect 2592 27716 2596 27772
rect 2596 27716 2652 27772
rect 2652 27716 2656 27772
rect 2592 27712 2656 27716
rect 33072 27772 33136 27776
rect 33072 27716 33076 27772
rect 33076 27716 33132 27772
rect 33132 27716 33136 27772
rect 33072 27712 33136 27716
rect 33152 27772 33216 27776
rect 33152 27716 33156 27772
rect 33156 27716 33212 27772
rect 33212 27716 33216 27772
rect 33152 27712 33216 27716
rect 33232 27772 33296 27776
rect 33232 27716 33236 27772
rect 33236 27716 33292 27772
rect 33292 27716 33296 27772
rect 33232 27712 33296 27716
rect 33312 27772 33376 27776
rect 33312 27716 33316 27772
rect 33316 27716 33372 27772
rect 33372 27716 33376 27772
rect 33312 27712 33376 27716
rect 3012 27228 3076 27232
rect 3012 27172 3016 27228
rect 3016 27172 3072 27228
rect 3072 27172 3076 27228
rect 3012 27168 3076 27172
rect 3092 27228 3156 27232
rect 3092 27172 3096 27228
rect 3096 27172 3152 27228
rect 3152 27172 3156 27228
rect 3092 27168 3156 27172
rect 3172 27228 3236 27232
rect 3172 27172 3176 27228
rect 3176 27172 3232 27228
rect 3232 27172 3236 27228
rect 3172 27168 3236 27172
rect 3252 27228 3316 27232
rect 3252 27172 3256 27228
rect 3256 27172 3312 27228
rect 3312 27172 3316 27228
rect 3252 27168 3316 27172
rect 33732 27228 33796 27232
rect 33732 27172 33736 27228
rect 33736 27172 33792 27228
rect 33792 27172 33796 27228
rect 33732 27168 33796 27172
rect 33812 27228 33876 27232
rect 33812 27172 33816 27228
rect 33816 27172 33872 27228
rect 33872 27172 33876 27228
rect 33812 27168 33876 27172
rect 33892 27228 33956 27232
rect 33892 27172 33896 27228
rect 33896 27172 33952 27228
rect 33952 27172 33956 27228
rect 33892 27168 33956 27172
rect 33972 27228 34036 27232
rect 33972 27172 33976 27228
rect 33976 27172 34032 27228
rect 34032 27172 34036 27228
rect 33972 27168 34036 27172
rect 2352 26684 2416 26688
rect 2352 26628 2356 26684
rect 2356 26628 2412 26684
rect 2412 26628 2416 26684
rect 2352 26624 2416 26628
rect 2432 26684 2496 26688
rect 2432 26628 2436 26684
rect 2436 26628 2492 26684
rect 2492 26628 2496 26684
rect 2432 26624 2496 26628
rect 2512 26684 2576 26688
rect 2512 26628 2516 26684
rect 2516 26628 2572 26684
rect 2572 26628 2576 26684
rect 2512 26624 2576 26628
rect 2592 26684 2656 26688
rect 2592 26628 2596 26684
rect 2596 26628 2652 26684
rect 2652 26628 2656 26684
rect 2592 26624 2656 26628
rect 33072 26684 33136 26688
rect 33072 26628 33076 26684
rect 33076 26628 33132 26684
rect 33132 26628 33136 26684
rect 33072 26624 33136 26628
rect 33152 26684 33216 26688
rect 33152 26628 33156 26684
rect 33156 26628 33212 26684
rect 33212 26628 33216 26684
rect 33152 26624 33216 26628
rect 33232 26684 33296 26688
rect 33232 26628 33236 26684
rect 33236 26628 33292 26684
rect 33292 26628 33296 26684
rect 33232 26624 33296 26628
rect 33312 26684 33376 26688
rect 33312 26628 33316 26684
rect 33316 26628 33372 26684
rect 33372 26628 33376 26684
rect 33312 26624 33376 26628
rect 3012 26140 3076 26144
rect 3012 26084 3016 26140
rect 3016 26084 3072 26140
rect 3072 26084 3076 26140
rect 3012 26080 3076 26084
rect 3092 26140 3156 26144
rect 3092 26084 3096 26140
rect 3096 26084 3152 26140
rect 3152 26084 3156 26140
rect 3092 26080 3156 26084
rect 3172 26140 3236 26144
rect 3172 26084 3176 26140
rect 3176 26084 3232 26140
rect 3232 26084 3236 26140
rect 3172 26080 3236 26084
rect 3252 26140 3316 26144
rect 3252 26084 3256 26140
rect 3256 26084 3312 26140
rect 3312 26084 3316 26140
rect 3252 26080 3316 26084
rect 33732 26140 33796 26144
rect 33732 26084 33736 26140
rect 33736 26084 33792 26140
rect 33792 26084 33796 26140
rect 33732 26080 33796 26084
rect 33812 26140 33876 26144
rect 33812 26084 33816 26140
rect 33816 26084 33872 26140
rect 33872 26084 33876 26140
rect 33812 26080 33876 26084
rect 33892 26140 33956 26144
rect 33892 26084 33896 26140
rect 33896 26084 33952 26140
rect 33952 26084 33956 26140
rect 33892 26080 33956 26084
rect 33972 26140 34036 26144
rect 33972 26084 33976 26140
rect 33976 26084 34032 26140
rect 34032 26084 34036 26140
rect 33972 26080 34036 26084
rect 2352 25596 2416 25600
rect 2352 25540 2356 25596
rect 2356 25540 2412 25596
rect 2412 25540 2416 25596
rect 2352 25536 2416 25540
rect 2432 25596 2496 25600
rect 2432 25540 2436 25596
rect 2436 25540 2492 25596
rect 2492 25540 2496 25596
rect 2432 25536 2496 25540
rect 2512 25596 2576 25600
rect 2512 25540 2516 25596
rect 2516 25540 2572 25596
rect 2572 25540 2576 25596
rect 2512 25536 2576 25540
rect 2592 25596 2656 25600
rect 2592 25540 2596 25596
rect 2596 25540 2652 25596
rect 2652 25540 2656 25596
rect 2592 25536 2656 25540
rect 33072 25596 33136 25600
rect 33072 25540 33076 25596
rect 33076 25540 33132 25596
rect 33132 25540 33136 25596
rect 33072 25536 33136 25540
rect 33152 25596 33216 25600
rect 33152 25540 33156 25596
rect 33156 25540 33212 25596
rect 33212 25540 33216 25596
rect 33152 25536 33216 25540
rect 33232 25596 33296 25600
rect 33232 25540 33236 25596
rect 33236 25540 33292 25596
rect 33292 25540 33296 25596
rect 33232 25536 33296 25540
rect 33312 25596 33376 25600
rect 33312 25540 33316 25596
rect 33316 25540 33372 25596
rect 33372 25540 33376 25596
rect 33312 25536 33376 25540
rect 3012 25052 3076 25056
rect 3012 24996 3016 25052
rect 3016 24996 3072 25052
rect 3072 24996 3076 25052
rect 3012 24992 3076 24996
rect 3092 25052 3156 25056
rect 3092 24996 3096 25052
rect 3096 24996 3152 25052
rect 3152 24996 3156 25052
rect 3092 24992 3156 24996
rect 3172 25052 3236 25056
rect 3172 24996 3176 25052
rect 3176 24996 3232 25052
rect 3232 24996 3236 25052
rect 3172 24992 3236 24996
rect 3252 25052 3316 25056
rect 3252 24996 3256 25052
rect 3256 24996 3312 25052
rect 3312 24996 3316 25052
rect 3252 24992 3316 24996
rect 33732 25052 33796 25056
rect 33732 24996 33736 25052
rect 33736 24996 33792 25052
rect 33792 24996 33796 25052
rect 33732 24992 33796 24996
rect 33812 25052 33876 25056
rect 33812 24996 33816 25052
rect 33816 24996 33872 25052
rect 33872 24996 33876 25052
rect 33812 24992 33876 24996
rect 33892 25052 33956 25056
rect 33892 24996 33896 25052
rect 33896 24996 33952 25052
rect 33952 24996 33956 25052
rect 33892 24992 33956 24996
rect 33972 25052 34036 25056
rect 33972 24996 33976 25052
rect 33976 24996 34032 25052
rect 34032 24996 34036 25052
rect 33972 24992 34036 24996
rect 2352 24508 2416 24512
rect 2352 24452 2356 24508
rect 2356 24452 2412 24508
rect 2412 24452 2416 24508
rect 2352 24448 2416 24452
rect 2432 24508 2496 24512
rect 2432 24452 2436 24508
rect 2436 24452 2492 24508
rect 2492 24452 2496 24508
rect 2432 24448 2496 24452
rect 2512 24508 2576 24512
rect 2512 24452 2516 24508
rect 2516 24452 2572 24508
rect 2572 24452 2576 24508
rect 2512 24448 2576 24452
rect 2592 24508 2656 24512
rect 2592 24452 2596 24508
rect 2596 24452 2652 24508
rect 2652 24452 2656 24508
rect 2592 24448 2656 24452
rect 33072 24508 33136 24512
rect 33072 24452 33076 24508
rect 33076 24452 33132 24508
rect 33132 24452 33136 24508
rect 33072 24448 33136 24452
rect 33152 24508 33216 24512
rect 33152 24452 33156 24508
rect 33156 24452 33212 24508
rect 33212 24452 33216 24508
rect 33152 24448 33216 24452
rect 33232 24508 33296 24512
rect 33232 24452 33236 24508
rect 33236 24452 33292 24508
rect 33292 24452 33296 24508
rect 33232 24448 33296 24452
rect 33312 24508 33376 24512
rect 33312 24452 33316 24508
rect 33316 24452 33372 24508
rect 33372 24452 33376 24508
rect 33312 24448 33376 24452
rect 3012 23964 3076 23968
rect 3012 23908 3016 23964
rect 3016 23908 3072 23964
rect 3072 23908 3076 23964
rect 3012 23904 3076 23908
rect 3092 23964 3156 23968
rect 3092 23908 3096 23964
rect 3096 23908 3152 23964
rect 3152 23908 3156 23964
rect 3092 23904 3156 23908
rect 3172 23964 3236 23968
rect 3172 23908 3176 23964
rect 3176 23908 3232 23964
rect 3232 23908 3236 23964
rect 3172 23904 3236 23908
rect 3252 23964 3316 23968
rect 3252 23908 3256 23964
rect 3256 23908 3312 23964
rect 3312 23908 3316 23964
rect 3252 23904 3316 23908
rect 33732 23964 33796 23968
rect 33732 23908 33736 23964
rect 33736 23908 33792 23964
rect 33792 23908 33796 23964
rect 33732 23904 33796 23908
rect 33812 23964 33876 23968
rect 33812 23908 33816 23964
rect 33816 23908 33872 23964
rect 33872 23908 33876 23964
rect 33812 23904 33876 23908
rect 33892 23964 33956 23968
rect 33892 23908 33896 23964
rect 33896 23908 33952 23964
rect 33952 23908 33956 23964
rect 33892 23904 33956 23908
rect 33972 23964 34036 23968
rect 33972 23908 33976 23964
rect 33976 23908 34032 23964
rect 34032 23908 34036 23964
rect 33972 23904 34036 23908
rect 2352 23420 2416 23424
rect 2352 23364 2356 23420
rect 2356 23364 2412 23420
rect 2412 23364 2416 23420
rect 2352 23360 2416 23364
rect 2432 23420 2496 23424
rect 2432 23364 2436 23420
rect 2436 23364 2492 23420
rect 2492 23364 2496 23420
rect 2432 23360 2496 23364
rect 2512 23420 2576 23424
rect 2512 23364 2516 23420
rect 2516 23364 2572 23420
rect 2572 23364 2576 23420
rect 2512 23360 2576 23364
rect 2592 23420 2656 23424
rect 2592 23364 2596 23420
rect 2596 23364 2652 23420
rect 2652 23364 2656 23420
rect 2592 23360 2656 23364
rect 33072 23420 33136 23424
rect 33072 23364 33076 23420
rect 33076 23364 33132 23420
rect 33132 23364 33136 23420
rect 33072 23360 33136 23364
rect 33152 23420 33216 23424
rect 33152 23364 33156 23420
rect 33156 23364 33212 23420
rect 33212 23364 33216 23420
rect 33152 23360 33216 23364
rect 33232 23420 33296 23424
rect 33232 23364 33236 23420
rect 33236 23364 33292 23420
rect 33292 23364 33296 23420
rect 33232 23360 33296 23364
rect 33312 23420 33376 23424
rect 33312 23364 33316 23420
rect 33316 23364 33372 23420
rect 33372 23364 33376 23420
rect 33312 23360 33376 23364
rect 3012 22876 3076 22880
rect 3012 22820 3016 22876
rect 3016 22820 3072 22876
rect 3072 22820 3076 22876
rect 3012 22816 3076 22820
rect 3092 22876 3156 22880
rect 3092 22820 3096 22876
rect 3096 22820 3152 22876
rect 3152 22820 3156 22876
rect 3092 22816 3156 22820
rect 3172 22876 3236 22880
rect 3172 22820 3176 22876
rect 3176 22820 3232 22876
rect 3232 22820 3236 22876
rect 3172 22816 3236 22820
rect 3252 22876 3316 22880
rect 3252 22820 3256 22876
rect 3256 22820 3312 22876
rect 3312 22820 3316 22876
rect 3252 22816 3316 22820
rect 33732 22876 33796 22880
rect 33732 22820 33736 22876
rect 33736 22820 33792 22876
rect 33792 22820 33796 22876
rect 33732 22816 33796 22820
rect 33812 22876 33876 22880
rect 33812 22820 33816 22876
rect 33816 22820 33872 22876
rect 33872 22820 33876 22876
rect 33812 22816 33876 22820
rect 33892 22876 33956 22880
rect 33892 22820 33896 22876
rect 33896 22820 33952 22876
rect 33952 22820 33956 22876
rect 33892 22816 33956 22820
rect 33972 22876 34036 22880
rect 33972 22820 33976 22876
rect 33976 22820 34032 22876
rect 34032 22820 34036 22876
rect 33972 22816 34036 22820
rect 2352 22332 2416 22336
rect 2352 22276 2356 22332
rect 2356 22276 2412 22332
rect 2412 22276 2416 22332
rect 2352 22272 2416 22276
rect 2432 22332 2496 22336
rect 2432 22276 2436 22332
rect 2436 22276 2492 22332
rect 2492 22276 2496 22332
rect 2432 22272 2496 22276
rect 2512 22332 2576 22336
rect 2512 22276 2516 22332
rect 2516 22276 2572 22332
rect 2572 22276 2576 22332
rect 2512 22272 2576 22276
rect 2592 22332 2656 22336
rect 2592 22276 2596 22332
rect 2596 22276 2652 22332
rect 2652 22276 2656 22332
rect 2592 22272 2656 22276
rect 33072 22332 33136 22336
rect 33072 22276 33076 22332
rect 33076 22276 33132 22332
rect 33132 22276 33136 22332
rect 33072 22272 33136 22276
rect 33152 22332 33216 22336
rect 33152 22276 33156 22332
rect 33156 22276 33212 22332
rect 33212 22276 33216 22332
rect 33152 22272 33216 22276
rect 33232 22332 33296 22336
rect 33232 22276 33236 22332
rect 33236 22276 33292 22332
rect 33292 22276 33296 22332
rect 33232 22272 33296 22276
rect 33312 22332 33376 22336
rect 33312 22276 33316 22332
rect 33316 22276 33372 22332
rect 33372 22276 33376 22332
rect 33312 22272 33376 22276
rect 3012 21788 3076 21792
rect 3012 21732 3016 21788
rect 3016 21732 3072 21788
rect 3072 21732 3076 21788
rect 3012 21728 3076 21732
rect 3092 21788 3156 21792
rect 3092 21732 3096 21788
rect 3096 21732 3152 21788
rect 3152 21732 3156 21788
rect 3092 21728 3156 21732
rect 3172 21788 3236 21792
rect 3172 21732 3176 21788
rect 3176 21732 3232 21788
rect 3232 21732 3236 21788
rect 3172 21728 3236 21732
rect 3252 21788 3316 21792
rect 3252 21732 3256 21788
rect 3256 21732 3312 21788
rect 3312 21732 3316 21788
rect 3252 21728 3316 21732
rect 33732 21788 33796 21792
rect 33732 21732 33736 21788
rect 33736 21732 33792 21788
rect 33792 21732 33796 21788
rect 33732 21728 33796 21732
rect 33812 21788 33876 21792
rect 33812 21732 33816 21788
rect 33816 21732 33872 21788
rect 33872 21732 33876 21788
rect 33812 21728 33876 21732
rect 33892 21788 33956 21792
rect 33892 21732 33896 21788
rect 33896 21732 33952 21788
rect 33952 21732 33956 21788
rect 33892 21728 33956 21732
rect 33972 21788 34036 21792
rect 33972 21732 33976 21788
rect 33976 21732 34032 21788
rect 34032 21732 34036 21788
rect 33972 21728 34036 21732
rect 2352 21244 2416 21248
rect 2352 21188 2356 21244
rect 2356 21188 2412 21244
rect 2412 21188 2416 21244
rect 2352 21184 2416 21188
rect 2432 21244 2496 21248
rect 2432 21188 2436 21244
rect 2436 21188 2492 21244
rect 2492 21188 2496 21244
rect 2432 21184 2496 21188
rect 2512 21244 2576 21248
rect 2512 21188 2516 21244
rect 2516 21188 2572 21244
rect 2572 21188 2576 21244
rect 2512 21184 2576 21188
rect 2592 21244 2656 21248
rect 2592 21188 2596 21244
rect 2596 21188 2652 21244
rect 2652 21188 2656 21244
rect 2592 21184 2656 21188
rect 33072 21244 33136 21248
rect 33072 21188 33076 21244
rect 33076 21188 33132 21244
rect 33132 21188 33136 21244
rect 33072 21184 33136 21188
rect 33152 21244 33216 21248
rect 33152 21188 33156 21244
rect 33156 21188 33212 21244
rect 33212 21188 33216 21244
rect 33152 21184 33216 21188
rect 33232 21244 33296 21248
rect 33232 21188 33236 21244
rect 33236 21188 33292 21244
rect 33292 21188 33296 21244
rect 33232 21184 33296 21188
rect 33312 21244 33376 21248
rect 33312 21188 33316 21244
rect 33316 21188 33372 21244
rect 33372 21188 33376 21244
rect 33312 21184 33376 21188
rect 3012 20700 3076 20704
rect 3012 20644 3016 20700
rect 3016 20644 3072 20700
rect 3072 20644 3076 20700
rect 3012 20640 3076 20644
rect 3092 20700 3156 20704
rect 3092 20644 3096 20700
rect 3096 20644 3152 20700
rect 3152 20644 3156 20700
rect 3092 20640 3156 20644
rect 3172 20700 3236 20704
rect 3172 20644 3176 20700
rect 3176 20644 3232 20700
rect 3232 20644 3236 20700
rect 3172 20640 3236 20644
rect 3252 20700 3316 20704
rect 3252 20644 3256 20700
rect 3256 20644 3312 20700
rect 3312 20644 3316 20700
rect 3252 20640 3316 20644
rect 33732 20700 33796 20704
rect 33732 20644 33736 20700
rect 33736 20644 33792 20700
rect 33792 20644 33796 20700
rect 33732 20640 33796 20644
rect 33812 20700 33876 20704
rect 33812 20644 33816 20700
rect 33816 20644 33872 20700
rect 33872 20644 33876 20700
rect 33812 20640 33876 20644
rect 33892 20700 33956 20704
rect 33892 20644 33896 20700
rect 33896 20644 33952 20700
rect 33952 20644 33956 20700
rect 33892 20640 33956 20644
rect 33972 20700 34036 20704
rect 33972 20644 33976 20700
rect 33976 20644 34032 20700
rect 34032 20644 34036 20700
rect 33972 20640 34036 20644
rect 2352 20156 2416 20160
rect 2352 20100 2356 20156
rect 2356 20100 2412 20156
rect 2412 20100 2416 20156
rect 2352 20096 2416 20100
rect 2432 20156 2496 20160
rect 2432 20100 2436 20156
rect 2436 20100 2492 20156
rect 2492 20100 2496 20156
rect 2432 20096 2496 20100
rect 2512 20156 2576 20160
rect 2512 20100 2516 20156
rect 2516 20100 2572 20156
rect 2572 20100 2576 20156
rect 2512 20096 2576 20100
rect 2592 20156 2656 20160
rect 2592 20100 2596 20156
rect 2596 20100 2652 20156
rect 2652 20100 2656 20156
rect 2592 20096 2656 20100
rect 33072 20156 33136 20160
rect 33072 20100 33076 20156
rect 33076 20100 33132 20156
rect 33132 20100 33136 20156
rect 33072 20096 33136 20100
rect 33152 20156 33216 20160
rect 33152 20100 33156 20156
rect 33156 20100 33212 20156
rect 33212 20100 33216 20156
rect 33152 20096 33216 20100
rect 33232 20156 33296 20160
rect 33232 20100 33236 20156
rect 33236 20100 33292 20156
rect 33292 20100 33296 20156
rect 33232 20096 33296 20100
rect 33312 20156 33376 20160
rect 33312 20100 33316 20156
rect 33316 20100 33372 20156
rect 33372 20100 33376 20156
rect 33312 20096 33376 20100
rect 3012 19612 3076 19616
rect 3012 19556 3016 19612
rect 3016 19556 3072 19612
rect 3072 19556 3076 19612
rect 3012 19552 3076 19556
rect 3092 19612 3156 19616
rect 3092 19556 3096 19612
rect 3096 19556 3152 19612
rect 3152 19556 3156 19612
rect 3092 19552 3156 19556
rect 3172 19612 3236 19616
rect 3172 19556 3176 19612
rect 3176 19556 3232 19612
rect 3232 19556 3236 19612
rect 3172 19552 3236 19556
rect 3252 19612 3316 19616
rect 3252 19556 3256 19612
rect 3256 19556 3312 19612
rect 3312 19556 3316 19612
rect 3252 19552 3316 19556
rect 33732 19612 33796 19616
rect 33732 19556 33736 19612
rect 33736 19556 33792 19612
rect 33792 19556 33796 19612
rect 33732 19552 33796 19556
rect 33812 19612 33876 19616
rect 33812 19556 33816 19612
rect 33816 19556 33872 19612
rect 33872 19556 33876 19612
rect 33812 19552 33876 19556
rect 33892 19612 33956 19616
rect 33892 19556 33896 19612
rect 33896 19556 33952 19612
rect 33952 19556 33956 19612
rect 33892 19552 33956 19556
rect 33972 19612 34036 19616
rect 33972 19556 33976 19612
rect 33976 19556 34032 19612
rect 34032 19556 34036 19612
rect 33972 19552 34036 19556
rect 2352 19068 2416 19072
rect 2352 19012 2356 19068
rect 2356 19012 2412 19068
rect 2412 19012 2416 19068
rect 2352 19008 2416 19012
rect 2432 19068 2496 19072
rect 2432 19012 2436 19068
rect 2436 19012 2492 19068
rect 2492 19012 2496 19068
rect 2432 19008 2496 19012
rect 2512 19068 2576 19072
rect 2512 19012 2516 19068
rect 2516 19012 2572 19068
rect 2572 19012 2576 19068
rect 2512 19008 2576 19012
rect 2592 19068 2656 19072
rect 2592 19012 2596 19068
rect 2596 19012 2652 19068
rect 2652 19012 2656 19068
rect 2592 19008 2656 19012
rect 33072 19068 33136 19072
rect 33072 19012 33076 19068
rect 33076 19012 33132 19068
rect 33132 19012 33136 19068
rect 33072 19008 33136 19012
rect 33152 19068 33216 19072
rect 33152 19012 33156 19068
rect 33156 19012 33212 19068
rect 33212 19012 33216 19068
rect 33152 19008 33216 19012
rect 33232 19068 33296 19072
rect 33232 19012 33236 19068
rect 33236 19012 33292 19068
rect 33292 19012 33296 19068
rect 33232 19008 33296 19012
rect 33312 19068 33376 19072
rect 33312 19012 33316 19068
rect 33316 19012 33372 19068
rect 33372 19012 33376 19068
rect 33312 19008 33376 19012
rect 3012 18524 3076 18528
rect 3012 18468 3016 18524
rect 3016 18468 3072 18524
rect 3072 18468 3076 18524
rect 3012 18464 3076 18468
rect 3092 18524 3156 18528
rect 3092 18468 3096 18524
rect 3096 18468 3152 18524
rect 3152 18468 3156 18524
rect 3092 18464 3156 18468
rect 3172 18524 3236 18528
rect 3172 18468 3176 18524
rect 3176 18468 3232 18524
rect 3232 18468 3236 18524
rect 3172 18464 3236 18468
rect 3252 18524 3316 18528
rect 3252 18468 3256 18524
rect 3256 18468 3312 18524
rect 3312 18468 3316 18524
rect 3252 18464 3316 18468
rect 33732 18524 33796 18528
rect 33732 18468 33736 18524
rect 33736 18468 33792 18524
rect 33792 18468 33796 18524
rect 33732 18464 33796 18468
rect 33812 18524 33876 18528
rect 33812 18468 33816 18524
rect 33816 18468 33872 18524
rect 33872 18468 33876 18524
rect 33812 18464 33876 18468
rect 33892 18524 33956 18528
rect 33892 18468 33896 18524
rect 33896 18468 33952 18524
rect 33952 18468 33956 18524
rect 33892 18464 33956 18468
rect 33972 18524 34036 18528
rect 33972 18468 33976 18524
rect 33976 18468 34032 18524
rect 34032 18468 34036 18524
rect 33972 18464 34036 18468
rect 2352 17980 2416 17984
rect 2352 17924 2356 17980
rect 2356 17924 2412 17980
rect 2412 17924 2416 17980
rect 2352 17920 2416 17924
rect 2432 17980 2496 17984
rect 2432 17924 2436 17980
rect 2436 17924 2492 17980
rect 2492 17924 2496 17980
rect 2432 17920 2496 17924
rect 2512 17980 2576 17984
rect 2512 17924 2516 17980
rect 2516 17924 2572 17980
rect 2572 17924 2576 17980
rect 2512 17920 2576 17924
rect 2592 17980 2656 17984
rect 2592 17924 2596 17980
rect 2596 17924 2652 17980
rect 2652 17924 2656 17980
rect 2592 17920 2656 17924
rect 33072 17980 33136 17984
rect 33072 17924 33076 17980
rect 33076 17924 33132 17980
rect 33132 17924 33136 17980
rect 33072 17920 33136 17924
rect 33152 17980 33216 17984
rect 33152 17924 33156 17980
rect 33156 17924 33212 17980
rect 33212 17924 33216 17980
rect 33152 17920 33216 17924
rect 33232 17980 33296 17984
rect 33232 17924 33236 17980
rect 33236 17924 33292 17980
rect 33292 17924 33296 17980
rect 33232 17920 33296 17924
rect 33312 17980 33376 17984
rect 33312 17924 33316 17980
rect 33316 17924 33372 17980
rect 33372 17924 33376 17980
rect 33312 17920 33376 17924
rect 3012 17436 3076 17440
rect 3012 17380 3016 17436
rect 3016 17380 3072 17436
rect 3072 17380 3076 17436
rect 3012 17376 3076 17380
rect 3092 17436 3156 17440
rect 3092 17380 3096 17436
rect 3096 17380 3152 17436
rect 3152 17380 3156 17436
rect 3092 17376 3156 17380
rect 3172 17436 3236 17440
rect 3172 17380 3176 17436
rect 3176 17380 3232 17436
rect 3232 17380 3236 17436
rect 3172 17376 3236 17380
rect 3252 17436 3316 17440
rect 3252 17380 3256 17436
rect 3256 17380 3312 17436
rect 3312 17380 3316 17436
rect 3252 17376 3316 17380
rect 33732 17436 33796 17440
rect 33732 17380 33736 17436
rect 33736 17380 33792 17436
rect 33792 17380 33796 17436
rect 33732 17376 33796 17380
rect 33812 17436 33876 17440
rect 33812 17380 33816 17436
rect 33816 17380 33872 17436
rect 33872 17380 33876 17436
rect 33812 17376 33876 17380
rect 33892 17436 33956 17440
rect 33892 17380 33896 17436
rect 33896 17380 33952 17436
rect 33952 17380 33956 17436
rect 33892 17376 33956 17380
rect 33972 17436 34036 17440
rect 33972 17380 33976 17436
rect 33976 17380 34032 17436
rect 34032 17380 34036 17436
rect 33972 17376 34036 17380
rect 2352 16892 2416 16896
rect 2352 16836 2356 16892
rect 2356 16836 2412 16892
rect 2412 16836 2416 16892
rect 2352 16832 2416 16836
rect 2432 16892 2496 16896
rect 2432 16836 2436 16892
rect 2436 16836 2492 16892
rect 2492 16836 2496 16892
rect 2432 16832 2496 16836
rect 2512 16892 2576 16896
rect 2512 16836 2516 16892
rect 2516 16836 2572 16892
rect 2572 16836 2576 16892
rect 2512 16832 2576 16836
rect 2592 16892 2656 16896
rect 2592 16836 2596 16892
rect 2596 16836 2652 16892
rect 2652 16836 2656 16892
rect 2592 16832 2656 16836
rect 33072 16892 33136 16896
rect 33072 16836 33076 16892
rect 33076 16836 33132 16892
rect 33132 16836 33136 16892
rect 33072 16832 33136 16836
rect 33152 16892 33216 16896
rect 33152 16836 33156 16892
rect 33156 16836 33212 16892
rect 33212 16836 33216 16892
rect 33152 16832 33216 16836
rect 33232 16892 33296 16896
rect 33232 16836 33236 16892
rect 33236 16836 33292 16892
rect 33292 16836 33296 16892
rect 33232 16832 33296 16836
rect 33312 16892 33376 16896
rect 33312 16836 33316 16892
rect 33316 16836 33372 16892
rect 33372 16836 33376 16892
rect 33312 16832 33376 16836
rect 3012 16348 3076 16352
rect 3012 16292 3016 16348
rect 3016 16292 3072 16348
rect 3072 16292 3076 16348
rect 3012 16288 3076 16292
rect 3092 16348 3156 16352
rect 3092 16292 3096 16348
rect 3096 16292 3152 16348
rect 3152 16292 3156 16348
rect 3092 16288 3156 16292
rect 3172 16348 3236 16352
rect 3172 16292 3176 16348
rect 3176 16292 3232 16348
rect 3232 16292 3236 16348
rect 3172 16288 3236 16292
rect 3252 16348 3316 16352
rect 3252 16292 3256 16348
rect 3256 16292 3312 16348
rect 3312 16292 3316 16348
rect 3252 16288 3316 16292
rect 33732 16348 33796 16352
rect 33732 16292 33736 16348
rect 33736 16292 33792 16348
rect 33792 16292 33796 16348
rect 33732 16288 33796 16292
rect 33812 16348 33876 16352
rect 33812 16292 33816 16348
rect 33816 16292 33872 16348
rect 33872 16292 33876 16348
rect 33812 16288 33876 16292
rect 33892 16348 33956 16352
rect 33892 16292 33896 16348
rect 33896 16292 33952 16348
rect 33952 16292 33956 16348
rect 33892 16288 33956 16292
rect 33972 16348 34036 16352
rect 33972 16292 33976 16348
rect 33976 16292 34032 16348
rect 34032 16292 34036 16348
rect 33972 16288 34036 16292
rect 2352 15804 2416 15808
rect 2352 15748 2356 15804
rect 2356 15748 2412 15804
rect 2412 15748 2416 15804
rect 2352 15744 2416 15748
rect 2432 15804 2496 15808
rect 2432 15748 2436 15804
rect 2436 15748 2492 15804
rect 2492 15748 2496 15804
rect 2432 15744 2496 15748
rect 2512 15804 2576 15808
rect 2512 15748 2516 15804
rect 2516 15748 2572 15804
rect 2572 15748 2576 15804
rect 2512 15744 2576 15748
rect 2592 15804 2656 15808
rect 2592 15748 2596 15804
rect 2596 15748 2652 15804
rect 2652 15748 2656 15804
rect 2592 15744 2656 15748
rect 33072 15804 33136 15808
rect 33072 15748 33076 15804
rect 33076 15748 33132 15804
rect 33132 15748 33136 15804
rect 33072 15744 33136 15748
rect 33152 15804 33216 15808
rect 33152 15748 33156 15804
rect 33156 15748 33212 15804
rect 33212 15748 33216 15804
rect 33152 15744 33216 15748
rect 33232 15804 33296 15808
rect 33232 15748 33236 15804
rect 33236 15748 33292 15804
rect 33292 15748 33296 15804
rect 33232 15744 33296 15748
rect 33312 15804 33376 15808
rect 33312 15748 33316 15804
rect 33316 15748 33372 15804
rect 33372 15748 33376 15804
rect 33312 15744 33376 15748
rect 3012 15260 3076 15264
rect 3012 15204 3016 15260
rect 3016 15204 3072 15260
rect 3072 15204 3076 15260
rect 3012 15200 3076 15204
rect 3092 15260 3156 15264
rect 3092 15204 3096 15260
rect 3096 15204 3152 15260
rect 3152 15204 3156 15260
rect 3092 15200 3156 15204
rect 3172 15260 3236 15264
rect 3172 15204 3176 15260
rect 3176 15204 3232 15260
rect 3232 15204 3236 15260
rect 3172 15200 3236 15204
rect 3252 15260 3316 15264
rect 3252 15204 3256 15260
rect 3256 15204 3312 15260
rect 3312 15204 3316 15260
rect 3252 15200 3316 15204
rect 33732 15260 33796 15264
rect 33732 15204 33736 15260
rect 33736 15204 33792 15260
rect 33792 15204 33796 15260
rect 33732 15200 33796 15204
rect 33812 15260 33876 15264
rect 33812 15204 33816 15260
rect 33816 15204 33872 15260
rect 33872 15204 33876 15260
rect 33812 15200 33876 15204
rect 33892 15260 33956 15264
rect 33892 15204 33896 15260
rect 33896 15204 33952 15260
rect 33952 15204 33956 15260
rect 33892 15200 33956 15204
rect 33972 15260 34036 15264
rect 33972 15204 33976 15260
rect 33976 15204 34032 15260
rect 34032 15204 34036 15260
rect 33972 15200 34036 15204
rect 2352 14716 2416 14720
rect 2352 14660 2356 14716
rect 2356 14660 2412 14716
rect 2412 14660 2416 14716
rect 2352 14656 2416 14660
rect 2432 14716 2496 14720
rect 2432 14660 2436 14716
rect 2436 14660 2492 14716
rect 2492 14660 2496 14716
rect 2432 14656 2496 14660
rect 2512 14716 2576 14720
rect 2512 14660 2516 14716
rect 2516 14660 2572 14716
rect 2572 14660 2576 14716
rect 2512 14656 2576 14660
rect 2592 14716 2656 14720
rect 2592 14660 2596 14716
rect 2596 14660 2652 14716
rect 2652 14660 2656 14716
rect 2592 14656 2656 14660
rect 33072 14716 33136 14720
rect 33072 14660 33076 14716
rect 33076 14660 33132 14716
rect 33132 14660 33136 14716
rect 33072 14656 33136 14660
rect 33152 14716 33216 14720
rect 33152 14660 33156 14716
rect 33156 14660 33212 14716
rect 33212 14660 33216 14716
rect 33152 14656 33216 14660
rect 33232 14716 33296 14720
rect 33232 14660 33236 14716
rect 33236 14660 33292 14716
rect 33292 14660 33296 14716
rect 33232 14656 33296 14660
rect 33312 14716 33376 14720
rect 33312 14660 33316 14716
rect 33316 14660 33372 14716
rect 33372 14660 33376 14716
rect 33312 14656 33376 14660
rect 3012 14172 3076 14176
rect 3012 14116 3016 14172
rect 3016 14116 3072 14172
rect 3072 14116 3076 14172
rect 3012 14112 3076 14116
rect 3092 14172 3156 14176
rect 3092 14116 3096 14172
rect 3096 14116 3152 14172
rect 3152 14116 3156 14172
rect 3092 14112 3156 14116
rect 3172 14172 3236 14176
rect 3172 14116 3176 14172
rect 3176 14116 3232 14172
rect 3232 14116 3236 14172
rect 3172 14112 3236 14116
rect 3252 14172 3316 14176
rect 3252 14116 3256 14172
rect 3256 14116 3312 14172
rect 3312 14116 3316 14172
rect 3252 14112 3316 14116
rect 33732 14172 33796 14176
rect 33732 14116 33736 14172
rect 33736 14116 33792 14172
rect 33792 14116 33796 14172
rect 33732 14112 33796 14116
rect 33812 14172 33876 14176
rect 33812 14116 33816 14172
rect 33816 14116 33872 14172
rect 33872 14116 33876 14172
rect 33812 14112 33876 14116
rect 33892 14172 33956 14176
rect 33892 14116 33896 14172
rect 33896 14116 33952 14172
rect 33952 14116 33956 14172
rect 33892 14112 33956 14116
rect 33972 14172 34036 14176
rect 33972 14116 33976 14172
rect 33976 14116 34032 14172
rect 34032 14116 34036 14172
rect 33972 14112 34036 14116
rect 2352 13628 2416 13632
rect 2352 13572 2356 13628
rect 2356 13572 2412 13628
rect 2412 13572 2416 13628
rect 2352 13568 2416 13572
rect 2432 13628 2496 13632
rect 2432 13572 2436 13628
rect 2436 13572 2492 13628
rect 2492 13572 2496 13628
rect 2432 13568 2496 13572
rect 2512 13628 2576 13632
rect 2512 13572 2516 13628
rect 2516 13572 2572 13628
rect 2572 13572 2576 13628
rect 2512 13568 2576 13572
rect 2592 13628 2656 13632
rect 2592 13572 2596 13628
rect 2596 13572 2652 13628
rect 2652 13572 2656 13628
rect 2592 13568 2656 13572
rect 33072 13628 33136 13632
rect 33072 13572 33076 13628
rect 33076 13572 33132 13628
rect 33132 13572 33136 13628
rect 33072 13568 33136 13572
rect 33152 13628 33216 13632
rect 33152 13572 33156 13628
rect 33156 13572 33212 13628
rect 33212 13572 33216 13628
rect 33152 13568 33216 13572
rect 33232 13628 33296 13632
rect 33232 13572 33236 13628
rect 33236 13572 33292 13628
rect 33292 13572 33296 13628
rect 33232 13568 33296 13572
rect 33312 13628 33376 13632
rect 33312 13572 33316 13628
rect 33316 13572 33372 13628
rect 33372 13572 33376 13628
rect 33312 13568 33376 13572
rect 3012 13084 3076 13088
rect 3012 13028 3016 13084
rect 3016 13028 3072 13084
rect 3072 13028 3076 13084
rect 3012 13024 3076 13028
rect 3092 13084 3156 13088
rect 3092 13028 3096 13084
rect 3096 13028 3152 13084
rect 3152 13028 3156 13084
rect 3092 13024 3156 13028
rect 3172 13084 3236 13088
rect 3172 13028 3176 13084
rect 3176 13028 3232 13084
rect 3232 13028 3236 13084
rect 3172 13024 3236 13028
rect 3252 13084 3316 13088
rect 3252 13028 3256 13084
rect 3256 13028 3312 13084
rect 3312 13028 3316 13084
rect 3252 13024 3316 13028
rect 33732 13084 33796 13088
rect 33732 13028 33736 13084
rect 33736 13028 33792 13084
rect 33792 13028 33796 13084
rect 33732 13024 33796 13028
rect 33812 13084 33876 13088
rect 33812 13028 33816 13084
rect 33816 13028 33872 13084
rect 33872 13028 33876 13084
rect 33812 13024 33876 13028
rect 33892 13084 33956 13088
rect 33892 13028 33896 13084
rect 33896 13028 33952 13084
rect 33952 13028 33956 13084
rect 33892 13024 33956 13028
rect 33972 13084 34036 13088
rect 33972 13028 33976 13084
rect 33976 13028 34032 13084
rect 34032 13028 34036 13084
rect 33972 13024 34036 13028
rect 2352 12540 2416 12544
rect 2352 12484 2356 12540
rect 2356 12484 2412 12540
rect 2412 12484 2416 12540
rect 2352 12480 2416 12484
rect 2432 12540 2496 12544
rect 2432 12484 2436 12540
rect 2436 12484 2492 12540
rect 2492 12484 2496 12540
rect 2432 12480 2496 12484
rect 2512 12540 2576 12544
rect 2512 12484 2516 12540
rect 2516 12484 2572 12540
rect 2572 12484 2576 12540
rect 2512 12480 2576 12484
rect 2592 12540 2656 12544
rect 2592 12484 2596 12540
rect 2596 12484 2652 12540
rect 2652 12484 2656 12540
rect 2592 12480 2656 12484
rect 33072 12540 33136 12544
rect 33072 12484 33076 12540
rect 33076 12484 33132 12540
rect 33132 12484 33136 12540
rect 33072 12480 33136 12484
rect 33152 12540 33216 12544
rect 33152 12484 33156 12540
rect 33156 12484 33212 12540
rect 33212 12484 33216 12540
rect 33152 12480 33216 12484
rect 33232 12540 33296 12544
rect 33232 12484 33236 12540
rect 33236 12484 33292 12540
rect 33292 12484 33296 12540
rect 33232 12480 33296 12484
rect 33312 12540 33376 12544
rect 33312 12484 33316 12540
rect 33316 12484 33372 12540
rect 33372 12484 33376 12540
rect 33312 12480 33376 12484
rect 3012 11996 3076 12000
rect 3012 11940 3016 11996
rect 3016 11940 3072 11996
rect 3072 11940 3076 11996
rect 3012 11936 3076 11940
rect 3092 11996 3156 12000
rect 3092 11940 3096 11996
rect 3096 11940 3152 11996
rect 3152 11940 3156 11996
rect 3092 11936 3156 11940
rect 3172 11996 3236 12000
rect 3172 11940 3176 11996
rect 3176 11940 3232 11996
rect 3232 11940 3236 11996
rect 3172 11936 3236 11940
rect 3252 11996 3316 12000
rect 3252 11940 3256 11996
rect 3256 11940 3312 11996
rect 3312 11940 3316 11996
rect 3252 11936 3316 11940
rect 33732 11996 33796 12000
rect 33732 11940 33736 11996
rect 33736 11940 33792 11996
rect 33792 11940 33796 11996
rect 33732 11936 33796 11940
rect 33812 11996 33876 12000
rect 33812 11940 33816 11996
rect 33816 11940 33872 11996
rect 33872 11940 33876 11996
rect 33812 11936 33876 11940
rect 33892 11996 33956 12000
rect 33892 11940 33896 11996
rect 33896 11940 33952 11996
rect 33952 11940 33956 11996
rect 33892 11936 33956 11940
rect 33972 11996 34036 12000
rect 33972 11940 33976 11996
rect 33976 11940 34032 11996
rect 34032 11940 34036 11996
rect 33972 11936 34036 11940
rect 2352 11452 2416 11456
rect 2352 11396 2356 11452
rect 2356 11396 2412 11452
rect 2412 11396 2416 11452
rect 2352 11392 2416 11396
rect 2432 11452 2496 11456
rect 2432 11396 2436 11452
rect 2436 11396 2492 11452
rect 2492 11396 2496 11452
rect 2432 11392 2496 11396
rect 2512 11452 2576 11456
rect 2512 11396 2516 11452
rect 2516 11396 2572 11452
rect 2572 11396 2576 11452
rect 2512 11392 2576 11396
rect 2592 11452 2656 11456
rect 2592 11396 2596 11452
rect 2596 11396 2652 11452
rect 2652 11396 2656 11452
rect 2592 11392 2656 11396
rect 33072 11452 33136 11456
rect 33072 11396 33076 11452
rect 33076 11396 33132 11452
rect 33132 11396 33136 11452
rect 33072 11392 33136 11396
rect 33152 11452 33216 11456
rect 33152 11396 33156 11452
rect 33156 11396 33212 11452
rect 33212 11396 33216 11452
rect 33152 11392 33216 11396
rect 33232 11452 33296 11456
rect 33232 11396 33236 11452
rect 33236 11396 33292 11452
rect 33292 11396 33296 11452
rect 33232 11392 33296 11396
rect 33312 11452 33376 11456
rect 33312 11396 33316 11452
rect 33316 11396 33372 11452
rect 33372 11396 33376 11452
rect 33312 11392 33376 11396
rect 3012 10908 3076 10912
rect 3012 10852 3016 10908
rect 3016 10852 3072 10908
rect 3072 10852 3076 10908
rect 3012 10848 3076 10852
rect 3092 10908 3156 10912
rect 3092 10852 3096 10908
rect 3096 10852 3152 10908
rect 3152 10852 3156 10908
rect 3092 10848 3156 10852
rect 3172 10908 3236 10912
rect 3172 10852 3176 10908
rect 3176 10852 3232 10908
rect 3232 10852 3236 10908
rect 3172 10848 3236 10852
rect 3252 10908 3316 10912
rect 3252 10852 3256 10908
rect 3256 10852 3312 10908
rect 3312 10852 3316 10908
rect 3252 10848 3316 10852
rect 33732 10908 33796 10912
rect 33732 10852 33736 10908
rect 33736 10852 33792 10908
rect 33792 10852 33796 10908
rect 33732 10848 33796 10852
rect 33812 10908 33876 10912
rect 33812 10852 33816 10908
rect 33816 10852 33872 10908
rect 33872 10852 33876 10908
rect 33812 10848 33876 10852
rect 33892 10908 33956 10912
rect 33892 10852 33896 10908
rect 33896 10852 33952 10908
rect 33952 10852 33956 10908
rect 33892 10848 33956 10852
rect 33972 10908 34036 10912
rect 33972 10852 33976 10908
rect 33976 10852 34032 10908
rect 34032 10852 34036 10908
rect 33972 10848 34036 10852
rect 2352 10364 2416 10368
rect 2352 10308 2356 10364
rect 2356 10308 2412 10364
rect 2412 10308 2416 10364
rect 2352 10304 2416 10308
rect 2432 10364 2496 10368
rect 2432 10308 2436 10364
rect 2436 10308 2492 10364
rect 2492 10308 2496 10364
rect 2432 10304 2496 10308
rect 2512 10364 2576 10368
rect 2512 10308 2516 10364
rect 2516 10308 2572 10364
rect 2572 10308 2576 10364
rect 2512 10304 2576 10308
rect 2592 10364 2656 10368
rect 2592 10308 2596 10364
rect 2596 10308 2652 10364
rect 2652 10308 2656 10364
rect 2592 10304 2656 10308
rect 33072 10364 33136 10368
rect 33072 10308 33076 10364
rect 33076 10308 33132 10364
rect 33132 10308 33136 10364
rect 33072 10304 33136 10308
rect 33152 10364 33216 10368
rect 33152 10308 33156 10364
rect 33156 10308 33212 10364
rect 33212 10308 33216 10364
rect 33152 10304 33216 10308
rect 33232 10364 33296 10368
rect 33232 10308 33236 10364
rect 33236 10308 33292 10364
rect 33292 10308 33296 10364
rect 33232 10304 33296 10308
rect 33312 10364 33376 10368
rect 33312 10308 33316 10364
rect 33316 10308 33372 10364
rect 33372 10308 33376 10364
rect 33312 10304 33376 10308
rect 3012 9820 3076 9824
rect 3012 9764 3016 9820
rect 3016 9764 3072 9820
rect 3072 9764 3076 9820
rect 3012 9760 3076 9764
rect 3092 9820 3156 9824
rect 3092 9764 3096 9820
rect 3096 9764 3152 9820
rect 3152 9764 3156 9820
rect 3092 9760 3156 9764
rect 3172 9820 3236 9824
rect 3172 9764 3176 9820
rect 3176 9764 3232 9820
rect 3232 9764 3236 9820
rect 3172 9760 3236 9764
rect 3252 9820 3316 9824
rect 3252 9764 3256 9820
rect 3256 9764 3312 9820
rect 3312 9764 3316 9820
rect 3252 9760 3316 9764
rect 33732 9820 33796 9824
rect 33732 9764 33736 9820
rect 33736 9764 33792 9820
rect 33792 9764 33796 9820
rect 33732 9760 33796 9764
rect 33812 9820 33876 9824
rect 33812 9764 33816 9820
rect 33816 9764 33872 9820
rect 33872 9764 33876 9820
rect 33812 9760 33876 9764
rect 33892 9820 33956 9824
rect 33892 9764 33896 9820
rect 33896 9764 33952 9820
rect 33952 9764 33956 9820
rect 33892 9760 33956 9764
rect 33972 9820 34036 9824
rect 33972 9764 33976 9820
rect 33976 9764 34032 9820
rect 34032 9764 34036 9820
rect 33972 9760 34036 9764
rect 2352 9276 2416 9280
rect 2352 9220 2356 9276
rect 2356 9220 2412 9276
rect 2412 9220 2416 9276
rect 2352 9216 2416 9220
rect 2432 9276 2496 9280
rect 2432 9220 2436 9276
rect 2436 9220 2492 9276
rect 2492 9220 2496 9276
rect 2432 9216 2496 9220
rect 2512 9276 2576 9280
rect 2512 9220 2516 9276
rect 2516 9220 2572 9276
rect 2572 9220 2576 9276
rect 2512 9216 2576 9220
rect 2592 9276 2656 9280
rect 2592 9220 2596 9276
rect 2596 9220 2652 9276
rect 2652 9220 2656 9276
rect 2592 9216 2656 9220
rect 33072 9276 33136 9280
rect 33072 9220 33076 9276
rect 33076 9220 33132 9276
rect 33132 9220 33136 9276
rect 33072 9216 33136 9220
rect 33152 9276 33216 9280
rect 33152 9220 33156 9276
rect 33156 9220 33212 9276
rect 33212 9220 33216 9276
rect 33152 9216 33216 9220
rect 33232 9276 33296 9280
rect 33232 9220 33236 9276
rect 33236 9220 33292 9276
rect 33292 9220 33296 9276
rect 33232 9216 33296 9220
rect 33312 9276 33376 9280
rect 33312 9220 33316 9276
rect 33316 9220 33372 9276
rect 33372 9220 33376 9276
rect 33312 9216 33376 9220
rect 3012 8732 3076 8736
rect 3012 8676 3016 8732
rect 3016 8676 3072 8732
rect 3072 8676 3076 8732
rect 3012 8672 3076 8676
rect 3092 8732 3156 8736
rect 3092 8676 3096 8732
rect 3096 8676 3152 8732
rect 3152 8676 3156 8732
rect 3092 8672 3156 8676
rect 3172 8732 3236 8736
rect 3172 8676 3176 8732
rect 3176 8676 3232 8732
rect 3232 8676 3236 8732
rect 3172 8672 3236 8676
rect 3252 8732 3316 8736
rect 3252 8676 3256 8732
rect 3256 8676 3312 8732
rect 3312 8676 3316 8732
rect 3252 8672 3316 8676
rect 33732 8732 33796 8736
rect 33732 8676 33736 8732
rect 33736 8676 33792 8732
rect 33792 8676 33796 8732
rect 33732 8672 33796 8676
rect 33812 8732 33876 8736
rect 33812 8676 33816 8732
rect 33816 8676 33872 8732
rect 33872 8676 33876 8732
rect 33812 8672 33876 8676
rect 33892 8732 33956 8736
rect 33892 8676 33896 8732
rect 33896 8676 33952 8732
rect 33952 8676 33956 8732
rect 33892 8672 33956 8676
rect 33972 8732 34036 8736
rect 33972 8676 33976 8732
rect 33976 8676 34032 8732
rect 34032 8676 34036 8732
rect 33972 8672 34036 8676
rect 2352 8188 2416 8192
rect 2352 8132 2356 8188
rect 2356 8132 2412 8188
rect 2412 8132 2416 8188
rect 2352 8128 2416 8132
rect 2432 8188 2496 8192
rect 2432 8132 2436 8188
rect 2436 8132 2492 8188
rect 2492 8132 2496 8188
rect 2432 8128 2496 8132
rect 2512 8188 2576 8192
rect 2512 8132 2516 8188
rect 2516 8132 2572 8188
rect 2572 8132 2576 8188
rect 2512 8128 2576 8132
rect 2592 8188 2656 8192
rect 2592 8132 2596 8188
rect 2596 8132 2652 8188
rect 2652 8132 2656 8188
rect 2592 8128 2656 8132
rect 33072 8188 33136 8192
rect 33072 8132 33076 8188
rect 33076 8132 33132 8188
rect 33132 8132 33136 8188
rect 33072 8128 33136 8132
rect 33152 8188 33216 8192
rect 33152 8132 33156 8188
rect 33156 8132 33212 8188
rect 33212 8132 33216 8188
rect 33152 8128 33216 8132
rect 33232 8188 33296 8192
rect 33232 8132 33236 8188
rect 33236 8132 33292 8188
rect 33292 8132 33296 8188
rect 33232 8128 33296 8132
rect 33312 8188 33376 8192
rect 33312 8132 33316 8188
rect 33316 8132 33372 8188
rect 33372 8132 33376 8188
rect 33312 8128 33376 8132
rect 3012 7644 3076 7648
rect 3012 7588 3016 7644
rect 3016 7588 3072 7644
rect 3072 7588 3076 7644
rect 3012 7584 3076 7588
rect 3092 7644 3156 7648
rect 3092 7588 3096 7644
rect 3096 7588 3152 7644
rect 3152 7588 3156 7644
rect 3092 7584 3156 7588
rect 3172 7644 3236 7648
rect 3172 7588 3176 7644
rect 3176 7588 3232 7644
rect 3232 7588 3236 7644
rect 3172 7584 3236 7588
rect 3252 7644 3316 7648
rect 3252 7588 3256 7644
rect 3256 7588 3312 7644
rect 3312 7588 3316 7644
rect 3252 7584 3316 7588
rect 33732 7644 33796 7648
rect 33732 7588 33736 7644
rect 33736 7588 33792 7644
rect 33792 7588 33796 7644
rect 33732 7584 33796 7588
rect 33812 7644 33876 7648
rect 33812 7588 33816 7644
rect 33816 7588 33872 7644
rect 33872 7588 33876 7644
rect 33812 7584 33876 7588
rect 33892 7644 33956 7648
rect 33892 7588 33896 7644
rect 33896 7588 33952 7644
rect 33952 7588 33956 7644
rect 33892 7584 33956 7588
rect 33972 7644 34036 7648
rect 33972 7588 33976 7644
rect 33976 7588 34032 7644
rect 34032 7588 34036 7644
rect 33972 7584 34036 7588
rect 2352 7100 2416 7104
rect 2352 7044 2356 7100
rect 2356 7044 2412 7100
rect 2412 7044 2416 7100
rect 2352 7040 2416 7044
rect 2432 7100 2496 7104
rect 2432 7044 2436 7100
rect 2436 7044 2492 7100
rect 2492 7044 2496 7100
rect 2432 7040 2496 7044
rect 2512 7100 2576 7104
rect 2512 7044 2516 7100
rect 2516 7044 2572 7100
rect 2572 7044 2576 7100
rect 2512 7040 2576 7044
rect 2592 7100 2656 7104
rect 2592 7044 2596 7100
rect 2596 7044 2652 7100
rect 2652 7044 2656 7100
rect 2592 7040 2656 7044
rect 33072 7100 33136 7104
rect 33072 7044 33076 7100
rect 33076 7044 33132 7100
rect 33132 7044 33136 7100
rect 33072 7040 33136 7044
rect 33152 7100 33216 7104
rect 33152 7044 33156 7100
rect 33156 7044 33212 7100
rect 33212 7044 33216 7100
rect 33152 7040 33216 7044
rect 33232 7100 33296 7104
rect 33232 7044 33236 7100
rect 33236 7044 33292 7100
rect 33292 7044 33296 7100
rect 33232 7040 33296 7044
rect 33312 7100 33376 7104
rect 33312 7044 33316 7100
rect 33316 7044 33372 7100
rect 33372 7044 33376 7100
rect 33312 7040 33376 7044
rect 3012 6556 3076 6560
rect 3012 6500 3016 6556
rect 3016 6500 3072 6556
rect 3072 6500 3076 6556
rect 3012 6496 3076 6500
rect 3092 6556 3156 6560
rect 3092 6500 3096 6556
rect 3096 6500 3152 6556
rect 3152 6500 3156 6556
rect 3092 6496 3156 6500
rect 3172 6556 3236 6560
rect 3172 6500 3176 6556
rect 3176 6500 3232 6556
rect 3232 6500 3236 6556
rect 3172 6496 3236 6500
rect 3252 6556 3316 6560
rect 3252 6500 3256 6556
rect 3256 6500 3312 6556
rect 3312 6500 3316 6556
rect 3252 6496 3316 6500
rect 33732 6556 33796 6560
rect 33732 6500 33736 6556
rect 33736 6500 33792 6556
rect 33792 6500 33796 6556
rect 33732 6496 33796 6500
rect 33812 6556 33876 6560
rect 33812 6500 33816 6556
rect 33816 6500 33872 6556
rect 33872 6500 33876 6556
rect 33812 6496 33876 6500
rect 33892 6556 33956 6560
rect 33892 6500 33896 6556
rect 33896 6500 33952 6556
rect 33952 6500 33956 6556
rect 33892 6496 33956 6500
rect 33972 6556 34036 6560
rect 33972 6500 33976 6556
rect 33976 6500 34032 6556
rect 34032 6500 34036 6556
rect 33972 6496 34036 6500
rect 2352 6012 2416 6016
rect 2352 5956 2356 6012
rect 2356 5956 2412 6012
rect 2412 5956 2416 6012
rect 2352 5952 2416 5956
rect 2432 6012 2496 6016
rect 2432 5956 2436 6012
rect 2436 5956 2492 6012
rect 2492 5956 2496 6012
rect 2432 5952 2496 5956
rect 2512 6012 2576 6016
rect 2512 5956 2516 6012
rect 2516 5956 2572 6012
rect 2572 5956 2576 6012
rect 2512 5952 2576 5956
rect 2592 6012 2656 6016
rect 2592 5956 2596 6012
rect 2596 5956 2652 6012
rect 2652 5956 2656 6012
rect 2592 5952 2656 5956
rect 33072 6012 33136 6016
rect 33072 5956 33076 6012
rect 33076 5956 33132 6012
rect 33132 5956 33136 6012
rect 33072 5952 33136 5956
rect 33152 6012 33216 6016
rect 33152 5956 33156 6012
rect 33156 5956 33212 6012
rect 33212 5956 33216 6012
rect 33152 5952 33216 5956
rect 33232 6012 33296 6016
rect 33232 5956 33236 6012
rect 33236 5956 33292 6012
rect 33292 5956 33296 6012
rect 33232 5952 33296 5956
rect 33312 6012 33376 6016
rect 33312 5956 33316 6012
rect 33316 5956 33372 6012
rect 33372 5956 33376 6012
rect 33312 5952 33376 5956
rect 3012 5468 3076 5472
rect 3012 5412 3016 5468
rect 3016 5412 3072 5468
rect 3072 5412 3076 5468
rect 3012 5408 3076 5412
rect 3092 5468 3156 5472
rect 3092 5412 3096 5468
rect 3096 5412 3152 5468
rect 3152 5412 3156 5468
rect 3092 5408 3156 5412
rect 3172 5468 3236 5472
rect 3172 5412 3176 5468
rect 3176 5412 3232 5468
rect 3232 5412 3236 5468
rect 3172 5408 3236 5412
rect 3252 5468 3316 5472
rect 3252 5412 3256 5468
rect 3256 5412 3312 5468
rect 3312 5412 3316 5468
rect 3252 5408 3316 5412
rect 33732 5468 33796 5472
rect 33732 5412 33736 5468
rect 33736 5412 33792 5468
rect 33792 5412 33796 5468
rect 33732 5408 33796 5412
rect 33812 5468 33876 5472
rect 33812 5412 33816 5468
rect 33816 5412 33872 5468
rect 33872 5412 33876 5468
rect 33812 5408 33876 5412
rect 33892 5468 33956 5472
rect 33892 5412 33896 5468
rect 33896 5412 33952 5468
rect 33952 5412 33956 5468
rect 33892 5408 33956 5412
rect 33972 5468 34036 5472
rect 33972 5412 33976 5468
rect 33976 5412 34032 5468
rect 34032 5412 34036 5468
rect 33972 5408 34036 5412
rect 2352 4924 2416 4928
rect 2352 4868 2356 4924
rect 2356 4868 2412 4924
rect 2412 4868 2416 4924
rect 2352 4864 2416 4868
rect 2432 4924 2496 4928
rect 2432 4868 2436 4924
rect 2436 4868 2492 4924
rect 2492 4868 2496 4924
rect 2432 4864 2496 4868
rect 2512 4924 2576 4928
rect 2512 4868 2516 4924
rect 2516 4868 2572 4924
rect 2572 4868 2576 4924
rect 2512 4864 2576 4868
rect 2592 4924 2656 4928
rect 2592 4868 2596 4924
rect 2596 4868 2652 4924
rect 2652 4868 2656 4924
rect 2592 4864 2656 4868
rect 33072 4924 33136 4928
rect 33072 4868 33076 4924
rect 33076 4868 33132 4924
rect 33132 4868 33136 4924
rect 33072 4864 33136 4868
rect 33152 4924 33216 4928
rect 33152 4868 33156 4924
rect 33156 4868 33212 4924
rect 33212 4868 33216 4924
rect 33152 4864 33216 4868
rect 33232 4924 33296 4928
rect 33232 4868 33236 4924
rect 33236 4868 33292 4924
rect 33292 4868 33296 4924
rect 33232 4864 33296 4868
rect 33312 4924 33376 4928
rect 33312 4868 33316 4924
rect 33316 4868 33372 4924
rect 33372 4868 33376 4924
rect 33312 4864 33376 4868
rect 3012 4380 3076 4384
rect 3012 4324 3016 4380
rect 3016 4324 3072 4380
rect 3072 4324 3076 4380
rect 3012 4320 3076 4324
rect 3092 4380 3156 4384
rect 3092 4324 3096 4380
rect 3096 4324 3152 4380
rect 3152 4324 3156 4380
rect 3092 4320 3156 4324
rect 3172 4380 3236 4384
rect 3172 4324 3176 4380
rect 3176 4324 3232 4380
rect 3232 4324 3236 4380
rect 3172 4320 3236 4324
rect 3252 4380 3316 4384
rect 3252 4324 3256 4380
rect 3256 4324 3312 4380
rect 3312 4324 3316 4380
rect 3252 4320 3316 4324
rect 33732 4380 33796 4384
rect 33732 4324 33736 4380
rect 33736 4324 33792 4380
rect 33792 4324 33796 4380
rect 33732 4320 33796 4324
rect 33812 4380 33876 4384
rect 33812 4324 33816 4380
rect 33816 4324 33872 4380
rect 33872 4324 33876 4380
rect 33812 4320 33876 4324
rect 33892 4380 33956 4384
rect 33892 4324 33896 4380
rect 33896 4324 33952 4380
rect 33952 4324 33956 4380
rect 33892 4320 33956 4324
rect 33972 4380 34036 4384
rect 33972 4324 33976 4380
rect 33976 4324 34032 4380
rect 34032 4324 34036 4380
rect 33972 4320 34036 4324
rect 2352 3836 2416 3840
rect 2352 3780 2356 3836
rect 2356 3780 2412 3836
rect 2412 3780 2416 3836
rect 2352 3776 2416 3780
rect 2432 3836 2496 3840
rect 2432 3780 2436 3836
rect 2436 3780 2492 3836
rect 2492 3780 2496 3836
rect 2432 3776 2496 3780
rect 2512 3836 2576 3840
rect 2512 3780 2516 3836
rect 2516 3780 2572 3836
rect 2572 3780 2576 3836
rect 2512 3776 2576 3780
rect 2592 3836 2656 3840
rect 2592 3780 2596 3836
rect 2596 3780 2652 3836
rect 2652 3780 2656 3836
rect 2592 3776 2656 3780
rect 33072 3836 33136 3840
rect 33072 3780 33076 3836
rect 33076 3780 33132 3836
rect 33132 3780 33136 3836
rect 33072 3776 33136 3780
rect 33152 3836 33216 3840
rect 33152 3780 33156 3836
rect 33156 3780 33212 3836
rect 33212 3780 33216 3836
rect 33152 3776 33216 3780
rect 33232 3836 33296 3840
rect 33232 3780 33236 3836
rect 33236 3780 33292 3836
rect 33292 3780 33296 3836
rect 33232 3776 33296 3780
rect 33312 3836 33376 3840
rect 33312 3780 33316 3836
rect 33316 3780 33372 3836
rect 33372 3780 33376 3836
rect 33312 3776 33376 3780
rect 3012 3292 3076 3296
rect 3012 3236 3016 3292
rect 3016 3236 3072 3292
rect 3072 3236 3076 3292
rect 3012 3232 3076 3236
rect 3092 3292 3156 3296
rect 3092 3236 3096 3292
rect 3096 3236 3152 3292
rect 3152 3236 3156 3292
rect 3092 3232 3156 3236
rect 3172 3292 3236 3296
rect 3172 3236 3176 3292
rect 3176 3236 3232 3292
rect 3232 3236 3236 3292
rect 3172 3232 3236 3236
rect 3252 3292 3316 3296
rect 3252 3236 3256 3292
rect 3256 3236 3312 3292
rect 3312 3236 3316 3292
rect 3252 3232 3316 3236
rect 33732 3292 33796 3296
rect 33732 3236 33736 3292
rect 33736 3236 33792 3292
rect 33792 3236 33796 3292
rect 33732 3232 33796 3236
rect 33812 3292 33876 3296
rect 33812 3236 33816 3292
rect 33816 3236 33872 3292
rect 33872 3236 33876 3292
rect 33812 3232 33876 3236
rect 33892 3292 33956 3296
rect 33892 3236 33896 3292
rect 33896 3236 33952 3292
rect 33952 3236 33956 3292
rect 33892 3232 33956 3236
rect 33972 3292 34036 3296
rect 33972 3236 33976 3292
rect 33976 3236 34032 3292
rect 34032 3236 34036 3292
rect 33972 3232 34036 3236
rect 2352 2748 2416 2752
rect 2352 2692 2356 2748
rect 2356 2692 2412 2748
rect 2412 2692 2416 2748
rect 2352 2688 2416 2692
rect 2432 2748 2496 2752
rect 2432 2692 2436 2748
rect 2436 2692 2492 2748
rect 2492 2692 2496 2748
rect 2432 2688 2496 2692
rect 2512 2748 2576 2752
rect 2512 2692 2516 2748
rect 2516 2692 2572 2748
rect 2572 2692 2576 2748
rect 2512 2688 2576 2692
rect 2592 2748 2656 2752
rect 2592 2692 2596 2748
rect 2596 2692 2652 2748
rect 2652 2692 2656 2748
rect 2592 2688 2656 2692
rect 33072 2748 33136 2752
rect 33072 2692 33076 2748
rect 33076 2692 33132 2748
rect 33132 2692 33136 2748
rect 33072 2688 33136 2692
rect 33152 2748 33216 2752
rect 33152 2692 33156 2748
rect 33156 2692 33212 2748
rect 33212 2692 33216 2748
rect 33152 2688 33216 2692
rect 33232 2748 33296 2752
rect 33232 2692 33236 2748
rect 33236 2692 33292 2748
rect 33292 2692 33296 2748
rect 33232 2688 33296 2692
rect 33312 2748 33376 2752
rect 33312 2692 33316 2748
rect 33316 2692 33372 2748
rect 33372 2692 33376 2748
rect 33312 2688 33376 2692
rect 3012 2204 3076 2208
rect 3012 2148 3016 2204
rect 3016 2148 3072 2204
rect 3072 2148 3076 2204
rect 3012 2144 3076 2148
rect 3092 2204 3156 2208
rect 3092 2148 3096 2204
rect 3096 2148 3152 2204
rect 3152 2148 3156 2204
rect 3092 2144 3156 2148
rect 3172 2204 3236 2208
rect 3172 2148 3176 2204
rect 3176 2148 3232 2204
rect 3232 2148 3236 2204
rect 3172 2144 3236 2148
rect 3252 2204 3316 2208
rect 3252 2148 3256 2204
rect 3256 2148 3312 2204
rect 3312 2148 3316 2204
rect 3252 2144 3316 2148
rect 33732 2204 33796 2208
rect 33732 2148 33736 2204
rect 33736 2148 33792 2204
rect 33792 2148 33796 2204
rect 33732 2144 33796 2148
rect 33812 2204 33876 2208
rect 33812 2148 33816 2204
rect 33816 2148 33872 2204
rect 33872 2148 33876 2204
rect 33812 2144 33876 2148
rect 33892 2204 33956 2208
rect 33892 2148 33896 2204
rect 33896 2148 33952 2204
rect 33952 2148 33956 2204
rect 33892 2144 33956 2148
rect 33972 2204 34036 2208
rect 33972 2148 33976 2204
rect 33976 2148 34032 2204
rect 34032 2148 34036 2204
rect 33972 2144 34036 2148
<< metal4 >>
rect 2344 57152 2664 57712
rect 2344 57088 2352 57152
rect 2416 57088 2432 57152
rect 2496 57088 2512 57152
rect 2576 57088 2592 57152
rect 2656 57088 2664 57152
rect 2344 56064 2664 57088
rect 2344 56000 2352 56064
rect 2416 56000 2432 56064
rect 2496 56000 2512 56064
rect 2576 56000 2592 56064
rect 2656 56000 2664 56064
rect 2344 54976 2664 56000
rect 2344 54912 2352 54976
rect 2416 54912 2432 54976
rect 2496 54912 2512 54976
rect 2576 54912 2592 54976
rect 2656 54912 2664 54976
rect 2344 53888 2664 54912
rect 2344 53824 2352 53888
rect 2416 53824 2432 53888
rect 2496 53824 2512 53888
rect 2576 53824 2592 53888
rect 2656 53824 2664 53888
rect 2344 52800 2664 53824
rect 2344 52736 2352 52800
rect 2416 52736 2432 52800
rect 2496 52736 2512 52800
rect 2576 52736 2592 52800
rect 2656 52736 2664 52800
rect 2344 51712 2664 52736
rect 2344 51648 2352 51712
rect 2416 51648 2432 51712
rect 2496 51648 2512 51712
rect 2576 51648 2592 51712
rect 2656 51648 2664 51712
rect 2344 50624 2664 51648
rect 2344 50560 2352 50624
rect 2416 50560 2432 50624
rect 2496 50560 2512 50624
rect 2576 50560 2592 50624
rect 2656 50560 2664 50624
rect 2344 49536 2664 50560
rect 2344 49472 2352 49536
rect 2416 49472 2432 49536
rect 2496 49472 2512 49536
rect 2576 49472 2592 49536
rect 2656 49472 2664 49536
rect 2344 48448 2664 49472
rect 2344 48384 2352 48448
rect 2416 48384 2432 48448
rect 2496 48384 2512 48448
rect 2576 48384 2592 48448
rect 2656 48384 2664 48448
rect 2344 47360 2664 48384
rect 2344 47296 2352 47360
rect 2416 47296 2432 47360
rect 2496 47296 2512 47360
rect 2576 47296 2592 47360
rect 2656 47296 2664 47360
rect 2344 46272 2664 47296
rect 2344 46208 2352 46272
rect 2416 46208 2432 46272
rect 2496 46208 2512 46272
rect 2576 46208 2592 46272
rect 2656 46208 2664 46272
rect 2344 45184 2664 46208
rect 2344 45120 2352 45184
rect 2416 45120 2432 45184
rect 2496 45120 2512 45184
rect 2576 45120 2592 45184
rect 2656 45120 2664 45184
rect 2344 44096 2664 45120
rect 2344 44032 2352 44096
rect 2416 44032 2432 44096
rect 2496 44032 2512 44096
rect 2576 44032 2592 44096
rect 2656 44032 2664 44096
rect 2344 43008 2664 44032
rect 2344 42944 2352 43008
rect 2416 42944 2432 43008
rect 2496 42944 2512 43008
rect 2576 42944 2592 43008
rect 2656 42944 2664 43008
rect 2344 41920 2664 42944
rect 2344 41856 2352 41920
rect 2416 41856 2432 41920
rect 2496 41856 2512 41920
rect 2576 41856 2592 41920
rect 2656 41856 2664 41920
rect 2344 40832 2664 41856
rect 2344 40768 2352 40832
rect 2416 40768 2432 40832
rect 2496 40768 2512 40832
rect 2576 40768 2592 40832
rect 2656 40768 2664 40832
rect 2344 39744 2664 40768
rect 2344 39680 2352 39744
rect 2416 39680 2432 39744
rect 2496 39680 2512 39744
rect 2576 39680 2592 39744
rect 2656 39680 2664 39744
rect 2344 38656 2664 39680
rect 2344 38592 2352 38656
rect 2416 38592 2432 38656
rect 2496 38592 2512 38656
rect 2576 38592 2592 38656
rect 2656 38592 2664 38656
rect 2344 37568 2664 38592
rect 2344 37504 2352 37568
rect 2416 37504 2432 37568
rect 2496 37504 2512 37568
rect 2576 37504 2592 37568
rect 2656 37504 2664 37568
rect 2344 36480 2664 37504
rect 2344 36416 2352 36480
rect 2416 36416 2432 36480
rect 2496 36416 2512 36480
rect 2576 36416 2592 36480
rect 2656 36416 2664 36480
rect 2344 35392 2664 36416
rect 2344 35328 2352 35392
rect 2416 35328 2432 35392
rect 2496 35328 2512 35392
rect 2576 35328 2592 35392
rect 2656 35328 2664 35392
rect 2344 34330 2664 35328
rect 2344 34304 2386 34330
rect 2622 34304 2664 34330
rect 2344 34240 2352 34304
rect 2656 34240 2664 34304
rect 2344 34094 2386 34240
rect 2622 34094 2664 34240
rect 2344 33216 2664 34094
rect 2344 33152 2352 33216
rect 2416 33152 2432 33216
rect 2496 33152 2512 33216
rect 2576 33152 2592 33216
rect 2656 33152 2664 33216
rect 2344 32128 2664 33152
rect 2344 32064 2352 32128
rect 2416 32064 2432 32128
rect 2496 32064 2512 32128
rect 2576 32064 2592 32128
rect 2656 32064 2664 32128
rect 2344 31040 2664 32064
rect 2344 30976 2352 31040
rect 2416 30976 2432 31040
rect 2496 30976 2512 31040
rect 2576 30976 2592 31040
rect 2656 30976 2664 31040
rect 2344 29952 2664 30976
rect 2344 29888 2352 29952
rect 2416 29888 2432 29952
rect 2496 29888 2512 29952
rect 2576 29888 2592 29952
rect 2656 29888 2664 29952
rect 2344 28864 2664 29888
rect 2344 28800 2352 28864
rect 2416 28800 2432 28864
rect 2496 28800 2512 28864
rect 2576 28800 2592 28864
rect 2656 28800 2664 28864
rect 2344 27776 2664 28800
rect 2344 27712 2352 27776
rect 2416 27712 2432 27776
rect 2496 27712 2512 27776
rect 2576 27712 2592 27776
rect 2656 27712 2664 27776
rect 2344 26688 2664 27712
rect 2344 26624 2352 26688
rect 2416 26624 2432 26688
rect 2496 26624 2512 26688
rect 2576 26624 2592 26688
rect 2656 26624 2664 26688
rect 2344 25600 2664 26624
rect 2344 25536 2352 25600
rect 2416 25536 2432 25600
rect 2496 25536 2512 25600
rect 2576 25536 2592 25600
rect 2656 25536 2664 25600
rect 2344 24512 2664 25536
rect 2344 24448 2352 24512
rect 2416 24448 2432 24512
rect 2496 24448 2512 24512
rect 2576 24448 2592 24512
rect 2656 24448 2664 24512
rect 2344 23424 2664 24448
rect 2344 23360 2352 23424
rect 2416 23360 2432 23424
rect 2496 23360 2512 23424
rect 2576 23360 2592 23424
rect 2656 23360 2664 23424
rect 2344 22336 2664 23360
rect 2344 22272 2352 22336
rect 2416 22272 2432 22336
rect 2496 22272 2512 22336
rect 2576 22272 2592 22336
rect 2656 22272 2664 22336
rect 2344 21248 2664 22272
rect 2344 21184 2352 21248
rect 2416 21184 2432 21248
rect 2496 21184 2512 21248
rect 2576 21184 2592 21248
rect 2656 21184 2664 21248
rect 2344 20160 2664 21184
rect 2344 20096 2352 20160
rect 2416 20096 2432 20160
rect 2496 20096 2512 20160
rect 2576 20096 2592 20160
rect 2656 20096 2664 20160
rect 2344 19072 2664 20096
rect 2344 19008 2352 19072
rect 2416 19008 2432 19072
rect 2496 19008 2512 19072
rect 2576 19008 2592 19072
rect 2656 19008 2664 19072
rect 2344 17984 2664 19008
rect 2344 17920 2352 17984
rect 2416 17920 2432 17984
rect 2496 17920 2512 17984
rect 2576 17920 2592 17984
rect 2656 17920 2664 17984
rect 2344 16896 2664 17920
rect 2344 16832 2352 16896
rect 2416 16832 2432 16896
rect 2496 16832 2512 16896
rect 2576 16832 2592 16896
rect 2656 16832 2664 16896
rect 2344 15808 2664 16832
rect 2344 15744 2352 15808
rect 2416 15744 2432 15808
rect 2496 15744 2512 15808
rect 2576 15744 2592 15808
rect 2656 15744 2664 15808
rect 2344 14720 2664 15744
rect 2344 14656 2352 14720
rect 2416 14656 2432 14720
rect 2496 14656 2512 14720
rect 2576 14656 2592 14720
rect 2656 14656 2664 14720
rect 2344 13632 2664 14656
rect 2344 13568 2352 13632
rect 2416 13568 2432 13632
rect 2496 13568 2512 13632
rect 2576 13568 2592 13632
rect 2656 13568 2664 13632
rect 2344 12544 2664 13568
rect 2344 12480 2352 12544
rect 2416 12480 2432 12544
rect 2496 12480 2512 12544
rect 2576 12480 2592 12544
rect 2656 12480 2664 12544
rect 2344 11456 2664 12480
rect 2344 11392 2352 11456
rect 2416 11392 2432 11456
rect 2496 11392 2512 11456
rect 2576 11392 2592 11456
rect 2656 11392 2664 11456
rect 2344 10368 2664 11392
rect 2344 10304 2352 10368
rect 2416 10304 2432 10368
rect 2496 10304 2512 10368
rect 2576 10304 2592 10368
rect 2656 10304 2664 10368
rect 2344 9280 2664 10304
rect 2344 9216 2352 9280
rect 2416 9216 2432 9280
rect 2496 9216 2512 9280
rect 2576 9216 2592 9280
rect 2656 9216 2664 9280
rect 2344 8192 2664 9216
rect 2344 8128 2352 8192
rect 2416 8128 2432 8192
rect 2496 8128 2512 8192
rect 2576 8128 2592 8192
rect 2656 8128 2664 8192
rect 2344 7104 2664 8128
rect 2344 7040 2352 7104
rect 2416 7040 2432 7104
rect 2496 7040 2512 7104
rect 2576 7040 2592 7104
rect 2656 7040 2664 7104
rect 2344 6016 2664 7040
rect 2344 5952 2352 6016
rect 2416 5952 2432 6016
rect 2496 5952 2512 6016
rect 2576 5952 2592 6016
rect 2656 5952 2664 6016
rect 2344 4928 2664 5952
rect 2344 4864 2352 4928
rect 2416 4864 2432 4928
rect 2496 4864 2512 4928
rect 2576 4864 2592 4928
rect 2656 4864 2664 4928
rect 2344 3840 2664 4864
rect 2344 3776 2352 3840
rect 2416 3776 2432 3840
rect 2496 3776 2512 3840
rect 2576 3776 2592 3840
rect 2656 3776 2664 3840
rect 2344 3694 2664 3776
rect 2344 3458 2386 3694
rect 2622 3458 2664 3694
rect 2344 2752 2664 3458
rect 2344 2688 2352 2752
rect 2416 2688 2432 2752
rect 2496 2688 2512 2752
rect 2576 2688 2592 2752
rect 2656 2688 2664 2752
rect 2344 2128 2664 2688
rect 3004 57696 3324 57712
rect 3004 57632 3012 57696
rect 3076 57632 3092 57696
rect 3156 57632 3172 57696
rect 3236 57632 3252 57696
rect 3316 57632 3324 57696
rect 3004 56608 3324 57632
rect 3004 56544 3012 56608
rect 3076 56544 3092 56608
rect 3156 56544 3172 56608
rect 3236 56544 3252 56608
rect 3316 56544 3324 56608
rect 3004 55520 3324 56544
rect 3004 55456 3012 55520
rect 3076 55456 3092 55520
rect 3156 55456 3172 55520
rect 3236 55456 3252 55520
rect 3316 55456 3324 55520
rect 3004 54432 3324 55456
rect 3004 54368 3012 54432
rect 3076 54368 3092 54432
rect 3156 54368 3172 54432
rect 3236 54368 3252 54432
rect 3316 54368 3324 54432
rect 3004 53344 3324 54368
rect 3004 53280 3012 53344
rect 3076 53280 3092 53344
rect 3156 53280 3172 53344
rect 3236 53280 3252 53344
rect 3316 53280 3324 53344
rect 3004 52256 3324 53280
rect 3004 52192 3012 52256
rect 3076 52192 3092 52256
rect 3156 52192 3172 52256
rect 3236 52192 3252 52256
rect 3316 52192 3324 52256
rect 3004 51168 3324 52192
rect 3004 51104 3012 51168
rect 3076 51104 3092 51168
rect 3156 51104 3172 51168
rect 3236 51104 3252 51168
rect 3316 51104 3324 51168
rect 3004 50080 3324 51104
rect 3004 50016 3012 50080
rect 3076 50016 3092 50080
rect 3156 50016 3172 50080
rect 3236 50016 3252 50080
rect 3316 50016 3324 50080
rect 3004 48992 3324 50016
rect 3004 48928 3012 48992
rect 3076 48928 3092 48992
rect 3156 48928 3172 48992
rect 3236 48928 3252 48992
rect 3316 48928 3324 48992
rect 3004 47904 3324 48928
rect 3004 47840 3012 47904
rect 3076 47840 3092 47904
rect 3156 47840 3172 47904
rect 3236 47840 3252 47904
rect 3316 47840 3324 47904
rect 3004 46816 3324 47840
rect 3004 46752 3012 46816
rect 3076 46752 3092 46816
rect 3156 46752 3172 46816
rect 3236 46752 3252 46816
rect 3316 46752 3324 46816
rect 3004 45728 3324 46752
rect 3004 45664 3012 45728
rect 3076 45664 3092 45728
rect 3156 45664 3172 45728
rect 3236 45664 3252 45728
rect 3316 45664 3324 45728
rect 3004 44640 3324 45664
rect 3004 44576 3012 44640
rect 3076 44576 3092 44640
rect 3156 44576 3172 44640
rect 3236 44576 3252 44640
rect 3316 44576 3324 44640
rect 3004 43552 3324 44576
rect 3004 43488 3012 43552
rect 3076 43488 3092 43552
rect 3156 43488 3172 43552
rect 3236 43488 3252 43552
rect 3316 43488 3324 43552
rect 3004 42464 3324 43488
rect 3004 42400 3012 42464
rect 3076 42400 3092 42464
rect 3156 42400 3172 42464
rect 3236 42400 3252 42464
rect 3316 42400 3324 42464
rect 3004 41376 3324 42400
rect 3004 41312 3012 41376
rect 3076 41312 3092 41376
rect 3156 41312 3172 41376
rect 3236 41312 3252 41376
rect 3316 41312 3324 41376
rect 3004 40288 3324 41312
rect 3004 40224 3012 40288
rect 3076 40224 3092 40288
rect 3156 40224 3172 40288
rect 3236 40224 3252 40288
rect 3316 40224 3324 40288
rect 3004 39200 3324 40224
rect 3004 39136 3012 39200
rect 3076 39136 3092 39200
rect 3156 39136 3172 39200
rect 3236 39136 3252 39200
rect 3316 39136 3324 39200
rect 3004 38112 3324 39136
rect 3004 38048 3012 38112
rect 3076 38048 3092 38112
rect 3156 38048 3172 38112
rect 3236 38048 3252 38112
rect 3316 38048 3324 38112
rect 3004 37024 3324 38048
rect 3004 36960 3012 37024
rect 3076 36960 3092 37024
rect 3156 36960 3172 37024
rect 3236 36960 3252 37024
rect 3316 36960 3324 37024
rect 3004 35936 3324 36960
rect 3004 35872 3012 35936
rect 3076 35872 3092 35936
rect 3156 35872 3172 35936
rect 3236 35872 3252 35936
rect 3316 35872 3324 35936
rect 3004 34990 3324 35872
rect 3004 34848 3046 34990
rect 3282 34848 3324 34990
rect 3004 34784 3012 34848
rect 3316 34784 3324 34848
rect 3004 34754 3046 34784
rect 3282 34754 3324 34784
rect 3004 33760 3324 34754
rect 3004 33696 3012 33760
rect 3076 33696 3092 33760
rect 3156 33696 3172 33760
rect 3236 33696 3252 33760
rect 3316 33696 3324 33760
rect 3004 32672 3324 33696
rect 3004 32608 3012 32672
rect 3076 32608 3092 32672
rect 3156 32608 3172 32672
rect 3236 32608 3252 32672
rect 3316 32608 3324 32672
rect 3004 31584 3324 32608
rect 3004 31520 3012 31584
rect 3076 31520 3092 31584
rect 3156 31520 3172 31584
rect 3236 31520 3252 31584
rect 3316 31520 3324 31584
rect 3004 30496 3324 31520
rect 3004 30432 3012 30496
rect 3076 30432 3092 30496
rect 3156 30432 3172 30496
rect 3236 30432 3252 30496
rect 3316 30432 3324 30496
rect 3004 29408 3324 30432
rect 3004 29344 3012 29408
rect 3076 29344 3092 29408
rect 3156 29344 3172 29408
rect 3236 29344 3252 29408
rect 3316 29344 3324 29408
rect 3004 28320 3324 29344
rect 3004 28256 3012 28320
rect 3076 28256 3092 28320
rect 3156 28256 3172 28320
rect 3236 28256 3252 28320
rect 3316 28256 3324 28320
rect 3004 27232 3324 28256
rect 3004 27168 3012 27232
rect 3076 27168 3092 27232
rect 3156 27168 3172 27232
rect 3236 27168 3252 27232
rect 3316 27168 3324 27232
rect 3004 26144 3324 27168
rect 3004 26080 3012 26144
rect 3076 26080 3092 26144
rect 3156 26080 3172 26144
rect 3236 26080 3252 26144
rect 3316 26080 3324 26144
rect 3004 25056 3324 26080
rect 3004 24992 3012 25056
rect 3076 24992 3092 25056
rect 3156 24992 3172 25056
rect 3236 24992 3252 25056
rect 3316 24992 3324 25056
rect 3004 23968 3324 24992
rect 3004 23904 3012 23968
rect 3076 23904 3092 23968
rect 3156 23904 3172 23968
rect 3236 23904 3252 23968
rect 3316 23904 3324 23968
rect 3004 22880 3324 23904
rect 3004 22816 3012 22880
rect 3076 22816 3092 22880
rect 3156 22816 3172 22880
rect 3236 22816 3252 22880
rect 3316 22816 3324 22880
rect 3004 21792 3324 22816
rect 3004 21728 3012 21792
rect 3076 21728 3092 21792
rect 3156 21728 3172 21792
rect 3236 21728 3252 21792
rect 3316 21728 3324 21792
rect 3004 20704 3324 21728
rect 3004 20640 3012 20704
rect 3076 20640 3092 20704
rect 3156 20640 3172 20704
rect 3236 20640 3252 20704
rect 3316 20640 3324 20704
rect 3004 19616 3324 20640
rect 3004 19552 3012 19616
rect 3076 19552 3092 19616
rect 3156 19552 3172 19616
rect 3236 19552 3252 19616
rect 3316 19552 3324 19616
rect 3004 18528 3324 19552
rect 3004 18464 3012 18528
rect 3076 18464 3092 18528
rect 3156 18464 3172 18528
rect 3236 18464 3252 18528
rect 3316 18464 3324 18528
rect 3004 17440 3324 18464
rect 3004 17376 3012 17440
rect 3076 17376 3092 17440
rect 3156 17376 3172 17440
rect 3236 17376 3252 17440
rect 3316 17376 3324 17440
rect 3004 16352 3324 17376
rect 3004 16288 3012 16352
rect 3076 16288 3092 16352
rect 3156 16288 3172 16352
rect 3236 16288 3252 16352
rect 3316 16288 3324 16352
rect 3004 15264 3324 16288
rect 3004 15200 3012 15264
rect 3076 15200 3092 15264
rect 3156 15200 3172 15264
rect 3236 15200 3252 15264
rect 3316 15200 3324 15264
rect 3004 14176 3324 15200
rect 3004 14112 3012 14176
rect 3076 14112 3092 14176
rect 3156 14112 3172 14176
rect 3236 14112 3252 14176
rect 3316 14112 3324 14176
rect 3004 13088 3324 14112
rect 3004 13024 3012 13088
rect 3076 13024 3092 13088
rect 3156 13024 3172 13088
rect 3236 13024 3252 13088
rect 3316 13024 3324 13088
rect 3004 12000 3324 13024
rect 3004 11936 3012 12000
rect 3076 11936 3092 12000
rect 3156 11936 3172 12000
rect 3236 11936 3252 12000
rect 3316 11936 3324 12000
rect 3004 10912 3324 11936
rect 3004 10848 3012 10912
rect 3076 10848 3092 10912
rect 3156 10848 3172 10912
rect 3236 10848 3252 10912
rect 3316 10848 3324 10912
rect 3004 9824 3324 10848
rect 3004 9760 3012 9824
rect 3076 9760 3092 9824
rect 3156 9760 3172 9824
rect 3236 9760 3252 9824
rect 3316 9760 3324 9824
rect 3004 8736 3324 9760
rect 3004 8672 3012 8736
rect 3076 8672 3092 8736
rect 3156 8672 3172 8736
rect 3236 8672 3252 8736
rect 3316 8672 3324 8736
rect 3004 7648 3324 8672
rect 3004 7584 3012 7648
rect 3076 7584 3092 7648
rect 3156 7584 3172 7648
rect 3236 7584 3252 7648
rect 3316 7584 3324 7648
rect 3004 6560 3324 7584
rect 3004 6496 3012 6560
rect 3076 6496 3092 6560
rect 3156 6496 3172 6560
rect 3236 6496 3252 6560
rect 3316 6496 3324 6560
rect 3004 5472 3324 6496
rect 3004 5408 3012 5472
rect 3076 5408 3092 5472
rect 3156 5408 3172 5472
rect 3236 5408 3252 5472
rect 3316 5408 3324 5472
rect 3004 4384 3324 5408
rect 3004 4320 3012 4384
rect 3076 4354 3092 4384
rect 3156 4354 3172 4384
rect 3236 4354 3252 4384
rect 3316 4320 3324 4384
rect 3004 4118 3046 4320
rect 3282 4118 3324 4320
rect 3004 3296 3324 4118
rect 3004 3232 3012 3296
rect 3076 3232 3092 3296
rect 3156 3232 3172 3296
rect 3236 3232 3252 3296
rect 3316 3232 3324 3296
rect 3004 2208 3324 3232
rect 3004 2144 3012 2208
rect 3076 2144 3092 2208
rect 3156 2144 3172 2208
rect 3236 2144 3252 2208
rect 3316 2144 3324 2208
rect 3004 2128 3324 2144
rect 33064 57152 33384 57712
rect 33064 57088 33072 57152
rect 33136 57088 33152 57152
rect 33216 57088 33232 57152
rect 33296 57088 33312 57152
rect 33376 57088 33384 57152
rect 33064 56064 33384 57088
rect 33064 56000 33072 56064
rect 33136 56000 33152 56064
rect 33216 56000 33232 56064
rect 33296 56000 33312 56064
rect 33376 56000 33384 56064
rect 33064 54976 33384 56000
rect 33064 54912 33072 54976
rect 33136 54912 33152 54976
rect 33216 54912 33232 54976
rect 33296 54912 33312 54976
rect 33376 54912 33384 54976
rect 33064 53888 33384 54912
rect 33064 53824 33072 53888
rect 33136 53824 33152 53888
rect 33216 53824 33232 53888
rect 33296 53824 33312 53888
rect 33376 53824 33384 53888
rect 33064 52800 33384 53824
rect 33064 52736 33072 52800
rect 33136 52736 33152 52800
rect 33216 52736 33232 52800
rect 33296 52736 33312 52800
rect 33376 52736 33384 52800
rect 33064 51712 33384 52736
rect 33064 51648 33072 51712
rect 33136 51648 33152 51712
rect 33216 51648 33232 51712
rect 33296 51648 33312 51712
rect 33376 51648 33384 51712
rect 33064 50624 33384 51648
rect 33064 50560 33072 50624
rect 33136 50560 33152 50624
rect 33216 50560 33232 50624
rect 33296 50560 33312 50624
rect 33376 50560 33384 50624
rect 33064 49536 33384 50560
rect 33064 49472 33072 49536
rect 33136 49472 33152 49536
rect 33216 49472 33232 49536
rect 33296 49472 33312 49536
rect 33376 49472 33384 49536
rect 33064 48448 33384 49472
rect 33064 48384 33072 48448
rect 33136 48384 33152 48448
rect 33216 48384 33232 48448
rect 33296 48384 33312 48448
rect 33376 48384 33384 48448
rect 33064 47360 33384 48384
rect 33064 47296 33072 47360
rect 33136 47296 33152 47360
rect 33216 47296 33232 47360
rect 33296 47296 33312 47360
rect 33376 47296 33384 47360
rect 33064 46272 33384 47296
rect 33064 46208 33072 46272
rect 33136 46208 33152 46272
rect 33216 46208 33232 46272
rect 33296 46208 33312 46272
rect 33376 46208 33384 46272
rect 33064 45184 33384 46208
rect 33064 45120 33072 45184
rect 33136 45120 33152 45184
rect 33216 45120 33232 45184
rect 33296 45120 33312 45184
rect 33376 45120 33384 45184
rect 33064 44096 33384 45120
rect 33064 44032 33072 44096
rect 33136 44032 33152 44096
rect 33216 44032 33232 44096
rect 33296 44032 33312 44096
rect 33376 44032 33384 44096
rect 33064 43008 33384 44032
rect 33064 42944 33072 43008
rect 33136 42944 33152 43008
rect 33216 42944 33232 43008
rect 33296 42944 33312 43008
rect 33376 42944 33384 43008
rect 33064 41920 33384 42944
rect 33064 41856 33072 41920
rect 33136 41856 33152 41920
rect 33216 41856 33232 41920
rect 33296 41856 33312 41920
rect 33376 41856 33384 41920
rect 33064 40832 33384 41856
rect 33064 40768 33072 40832
rect 33136 40768 33152 40832
rect 33216 40768 33232 40832
rect 33296 40768 33312 40832
rect 33376 40768 33384 40832
rect 33064 39744 33384 40768
rect 33064 39680 33072 39744
rect 33136 39680 33152 39744
rect 33216 39680 33232 39744
rect 33296 39680 33312 39744
rect 33376 39680 33384 39744
rect 33064 38656 33384 39680
rect 33064 38592 33072 38656
rect 33136 38592 33152 38656
rect 33216 38592 33232 38656
rect 33296 38592 33312 38656
rect 33376 38592 33384 38656
rect 33064 37568 33384 38592
rect 33064 37504 33072 37568
rect 33136 37504 33152 37568
rect 33216 37504 33232 37568
rect 33296 37504 33312 37568
rect 33376 37504 33384 37568
rect 33064 36480 33384 37504
rect 33064 36416 33072 36480
rect 33136 36416 33152 36480
rect 33216 36416 33232 36480
rect 33296 36416 33312 36480
rect 33376 36416 33384 36480
rect 33064 35392 33384 36416
rect 33064 35328 33072 35392
rect 33136 35328 33152 35392
rect 33216 35328 33232 35392
rect 33296 35328 33312 35392
rect 33376 35328 33384 35392
rect 33064 34330 33384 35328
rect 33064 34304 33106 34330
rect 33342 34304 33384 34330
rect 33064 34240 33072 34304
rect 33376 34240 33384 34304
rect 33064 34094 33106 34240
rect 33342 34094 33384 34240
rect 33064 33216 33384 34094
rect 33064 33152 33072 33216
rect 33136 33152 33152 33216
rect 33216 33152 33232 33216
rect 33296 33152 33312 33216
rect 33376 33152 33384 33216
rect 33064 32128 33384 33152
rect 33064 32064 33072 32128
rect 33136 32064 33152 32128
rect 33216 32064 33232 32128
rect 33296 32064 33312 32128
rect 33376 32064 33384 32128
rect 33064 31040 33384 32064
rect 33064 30976 33072 31040
rect 33136 30976 33152 31040
rect 33216 30976 33232 31040
rect 33296 30976 33312 31040
rect 33376 30976 33384 31040
rect 33064 29952 33384 30976
rect 33064 29888 33072 29952
rect 33136 29888 33152 29952
rect 33216 29888 33232 29952
rect 33296 29888 33312 29952
rect 33376 29888 33384 29952
rect 33064 28864 33384 29888
rect 33064 28800 33072 28864
rect 33136 28800 33152 28864
rect 33216 28800 33232 28864
rect 33296 28800 33312 28864
rect 33376 28800 33384 28864
rect 33064 27776 33384 28800
rect 33064 27712 33072 27776
rect 33136 27712 33152 27776
rect 33216 27712 33232 27776
rect 33296 27712 33312 27776
rect 33376 27712 33384 27776
rect 33064 26688 33384 27712
rect 33064 26624 33072 26688
rect 33136 26624 33152 26688
rect 33216 26624 33232 26688
rect 33296 26624 33312 26688
rect 33376 26624 33384 26688
rect 33064 25600 33384 26624
rect 33064 25536 33072 25600
rect 33136 25536 33152 25600
rect 33216 25536 33232 25600
rect 33296 25536 33312 25600
rect 33376 25536 33384 25600
rect 33064 24512 33384 25536
rect 33064 24448 33072 24512
rect 33136 24448 33152 24512
rect 33216 24448 33232 24512
rect 33296 24448 33312 24512
rect 33376 24448 33384 24512
rect 33064 23424 33384 24448
rect 33064 23360 33072 23424
rect 33136 23360 33152 23424
rect 33216 23360 33232 23424
rect 33296 23360 33312 23424
rect 33376 23360 33384 23424
rect 33064 22336 33384 23360
rect 33064 22272 33072 22336
rect 33136 22272 33152 22336
rect 33216 22272 33232 22336
rect 33296 22272 33312 22336
rect 33376 22272 33384 22336
rect 33064 21248 33384 22272
rect 33064 21184 33072 21248
rect 33136 21184 33152 21248
rect 33216 21184 33232 21248
rect 33296 21184 33312 21248
rect 33376 21184 33384 21248
rect 33064 20160 33384 21184
rect 33064 20096 33072 20160
rect 33136 20096 33152 20160
rect 33216 20096 33232 20160
rect 33296 20096 33312 20160
rect 33376 20096 33384 20160
rect 33064 19072 33384 20096
rect 33064 19008 33072 19072
rect 33136 19008 33152 19072
rect 33216 19008 33232 19072
rect 33296 19008 33312 19072
rect 33376 19008 33384 19072
rect 33064 17984 33384 19008
rect 33064 17920 33072 17984
rect 33136 17920 33152 17984
rect 33216 17920 33232 17984
rect 33296 17920 33312 17984
rect 33376 17920 33384 17984
rect 33064 16896 33384 17920
rect 33064 16832 33072 16896
rect 33136 16832 33152 16896
rect 33216 16832 33232 16896
rect 33296 16832 33312 16896
rect 33376 16832 33384 16896
rect 33064 15808 33384 16832
rect 33064 15744 33072 15808
rect 33136 15744 33152 15808
rect 33216 15744 33232 15808
rect 33296 15744 33312 15808
rect 33376 15744 33384 15808
rect 33064 14720 33384 15744
rect 33064 14656 33072 14720
rect 33136 14656 33152 14720
rect 33216 14656 33232 14720
rect 33296 14656 33312 14720
rect 33376 14656 33384 14720
rect 33064 13632 33384 14656
rect 33064 13568 33072 13632
rect 33136 13568 33152 13632
rect 33216 13568 33232 13632
rect 33296 13568 33312 13632
rect 33376 13568 33384 13632
rect 33064 12544 33384 13568
rect 33064 12480 33072 12544
rect 33136 12480 33152 12544
rect 33216 12480 33232 12544
rect 33296 12480 33312 12544
rect 33376 12480 33384 12544
rect 33064 11456 33384 12480
rect 33064 11392 33072 11456
rect 33136 11392 33152 11456
rect 33216 11392 33232 11456
rect 33296 11392 33312 11456
rect 33376 11392 33384 11456
rect 33064 10368 33384 11392
rect 33064 10304 33072 10368
rect 33136 10304 33152 10368
rect 33216 10304 33232 10368
rect 33296 10304 33312 10368
rect 33376 10304 33384 10368
rect 33064 9280 33384 10304
rect 33064 9216 33072 9280
rect 33136 9216 33152 9280
rect 33216 9216 33232 9280
rect 33296 9216 33312 9280
rect 33376 9216 33384 9280
rect 33064 8192 33384 9216
rect 33064 8128 33072 8192
rect 33136 8128 33152 8192
rect 33216 8128 33232 8192
rect 33296 8128 33312 8192
rect 33376 8128 33384 8192
rect 33064 7104 33384 8128
rect 33064 7040 33072 7104
rect 33136 7040 33152 7104
rect 33216 7040 33232 7104
rect 33296 7040 33312 7104
rect 33376 7040 33384 7104
rect 33064 6016 33384 7040
rect 33064 5952 33072 6016
rect 33136 5952 33152 6016
rect 33216 5952 33232 6016
rect 33296 5952 33312 6016
rect 33376 5952 33384 6016
rect 33064 4928 33384 5952
rect 33064 4864 33072 4928
rect 33136 4864 33152 4928
rect 33216 4864 33232 4928
rect 33296 4864 33312 4928
rect 33376 4864 33384 4928
rect 33064 3840 33384 4864
rect 33064 3776 33072 3840
rect 33136 3776 33152 3840
rect 33216 3776 33232 3840
rect 33296 3776 33312 3840
rect 33376 3776 33384 3840
rect 33064 3694 33384 3776
rect 33064 3458 33106 3694
rect 33342 3458 33384 3694
rect 33064 2752 33384 3458
rect 33064 2688 33072 2752
rect 33136 2688 33152 2752
rect 33216 2688 33232 2752
rect 33296 2688 33312 2752
rect 33376 2688 33384 2752
rect 33064 2128 33384 2688
rect 33724 57696 34044 57712
rect 33724 57632 33732 57696
rect 33796 57632 33812 57696
rect 33876 57632 33892 57696
rect 33956 57632 33972 57696
rect 34036 57632 34044 57696
rect 33724 56608 34044 57632
rect 33724 56544 33732 56608
rect 33796 56544 33812 56608
rect 33876 56544 33892 56608
rect 33956 56544 33972 56608
rect 34036 56544 34044 56608
rect 33724 55520 34044 56544
rect 33724 55456 33732 55520
rect 33796 55456 33812 55520
rect 33876 55456 33892 55520
rect 33956 55456 33972 55520
rect 34036 55456 34044 55520
rect 33724 54432 34044 55456
rect 33724 54368 33732 54432
rect 33796 54368 33812 54432
rect 33876 54368 33892 54432
rect 33956 54368 33972 54432
rect 34036 54368 34044 54432
rect 33724 53344 34044 54368
rect 33724 53280 33732 53344
rect 33796 53280 33812 53344
rect 33876 53280 33892 53344
rect 33956 53280 33972 53344
rect 34036 53280 34044 53344
rect 33724 52256 34044 53280
rect 33724 52192 33732 52256
rect 33796 52192 33812 52256
rect 33876 52192 33892 52256
rect 33956 52192 33972 52256
rect 34036 52192 34044 52256
rect 33724 51168 34044 52192
rect 33724 51104 33732 51168
rect 33796 51104 33812 51168
rect 33876 51104 33892 51168
rect 33956 51104 33972 51168
rect 34036 51104 34044 51168
rect 33724 50080 34044 51104
rect 33724 50016 33732 50080
rect 33796 50016 33812 50080
rect 33876 50016 33892 50080
rect 33956 50016 33972 50080
rect 34036 50016 34044 50080
rect 33724 48992 34044 50016
rect 33724 48928 33732 48992
rect 33796 48928 33812 48992
rect 33876 48928 33892 48992
rect 33956 48928 33972 48992
rect 34036 48928 34044 48992
rect 33724 47904 34044 48928
rect 33724 47840 33732 47904
rect 33796 47840 33812 47904
rect 33876 47840 33892 47904
rect 33956 47840 33972 47904
rect 34036 47840 34044 47904
rect 33724 46816 34044 47840
rect 33724 46752 33732 46816
rect 33796 46752 33812 46816
rect 33876 46752 33892 46816
rect 33956 46752 33972 46816
rect 34036 46752 34044 46816
rect 33724 45728 34044 46752
rect 33724 45664 33732 45728
rect 33796 45664 33812 45728
rect 33876 45664 33892 45728
rect 33956 45664 33972 45728
rect 34036 45664 34044 45728
rect 33724 44640 34044 45664
rect 33724 44576 33732 44640
rect 33796 44576 33812 44640
rect 33876 44576 33892 44640
rect 33956 44576 33972 44640
rect 34036 44576 34044 44640
rect 33724 43552 34044 44576
rect 33724 43488 33732 43552
rect 33796 43488 33812 43552
rect 33876 43488 33892 43552
rect 33956 43488 33972 43552
rect 34036 43488 34044 43552
rect 33724 42464 34044 43488
rect 33724 42400 33732 42464
rect 33796 42400 33812 42464
rect 33876 42400 33892 42464
rect 33956 42400 33972 42464
rect 34036 42400 34044 42464
rect 33724 41376 34044 42400
rect 33724 41312 33732 41376
rect 33796 41312 33812 41376
rect 33876 41312 33892 41376
rect 33956 41312 33972 41376
rect 34036 41312 34044 41376
rect 33724 40288 34044 41312
rect 33724 40224 33732 40288
rect 33796 40224 33812 40288
rect 33876 40224 33892 40288
rect 33956 40224 33972 40288
rect 34036 40224 34044 40288
rect 33724 39200 34044 40224
rect 33724 39136 33732 39200
rect 33796 39136 33812 39200
rect 33876 39136 33892 39200
rect 33956 39136 33972 39200
rect 34036 39136 34044 39200
rect 33724 38112 34044 39136
rect 33724 38048 33732 38112
rect 33796 38048 33812 38112
rect 33876 38048 33892 38112
rect 33956 38048 33972 38112
rect 34036 38048 34044 38112
rect 33724 37024 34044 38048
rect 33724 36960 33732 37024
rect 33796 36960 33812 37024
rect 33876 36960 33892 37024
rect 33956 36960 33972 37024
rect 34036 36960 34044 37024
rect 33724 35936 34044 36960
rect 33724 35872 33732 35936
rect 33796 35872 33812 35936
rect 33876 35872 33892 35936
rect 33956 35872 33972 35936
rect 34036 35872 34044 35936
rect 33724 34990 34044 35872
rect 33724 34848 33766 34990
rect 34002 34848 34044 34990
rect 33724 34784 33732 34848
rect 34036 34784 34044 34848
rect 33724 34754 33766 34784
rect 34002 34754 34044 34784
rect 33724 33760 34044 34754
rect 33724 33696 33732 33760
rect 33796 33696 33812 33760
rect 33876 33696 33892 33760
rect 33956 33696 33972 33760
rect 34036 33696 34044 33760
rect 33724 32672 34044 33696
rect 33724 32608 33732 32672
rect 33796 32608 33812 32672
rect 33876 32608 33892 32672
rect 33956 32608 33972 32672
rect 34036 32608 34044 32672
rect 33724 31584 34044 32608
rect 33724 31520 33732 31584
rect 33796 31520 33812 31584
rect 33876 31520 33892 31584
rect 33956 31520 33972 31584
rect 34036 31520 34044 31584
rect 33724 30496 34044 31520
rect 33724 30432 33732 30496
rect 33796 30432 33812 30496
rect 33876 30432 33892 30496
rect 33956 30432 33972 30496
rect 34036 30432 34044 30496
rect 33724 29408 34044 30432
rect 33724 29344 33732 29408
rect 33796 29344 33812 29408
rect 33876 29344 33892 29408
rect 33956 29344 33972 29408
rect 34036 29344 34044 29408
rect 33724 28320 34044 29344
rect 33724 28256 33732 28320
rect 33796 28256 33812 28320
rect 33876 28256 33892 28320
rect 33956 28256 33972 28320
rect 34036 28256 34044 28320
rect 33724 27232 34044 28256
rect 33724 27168 33732 27232
rect 33796 27168 33812 27232
rect 33876 27168 33892 27232
rect 33956 27168 33972 27232
rect 34036 27168 34044 27232
rect 33724 26144 34044 27168
rect 33724 26080 33732 26144
rect 33796 26080 33812 26144
rect 33876 26080 33892 26144
rect 33956 26080 33972 26144
rect 34036 26080 34044 26144
rect 33724 25056 34044 26080
rect 33724 24992 33732 25056
rect 33796 24992 33812 25056
rect 33876 24992 33892 25056
rect 33956 24992 33972 25056
rect 34036 24992 34044 25056
rect 33724 23968 34044 24992
rect 33724 23904 33732 23968
rect 33796 23904 33812 23968
rect 33876 23904 33892 23968
rect 33956 23904 33972 23968
rect 34036 23904 34044 23968
rect 33724 22880 34044 23904
rect 33724 22816 33732 22880
rect 33796 22816 33812 22880
rect 33876 22816 33892 22880
rect 33956 22816 33972 22880
rect 34036 22816 34044 22880
rect 33724 21792 34044 22816
rect 33724 21728 33732 21792
rect 33796 21728 33812 21792
rect 33876 21728 33892 21792
rect 33956 21728 33972 21792
rect 34036 21728 34044 21792
rect 33724 20704 34044 21728
rect 33724 20640 33732 20704
rect 33796 20640 33812 20704
rect 33876 20640 33892 20704
rect 33956 20640 33972 20704
rect 34036 20640 34044 20704
rect 33724 19616 34044 20640
rect 33724 19552 33732 19616
rect 33796 19552 33812 19616
rect 33876 19552 33892 19616
rect 33956 19552 33972 19616
rect 34036 19552 34044 19616
rect 33724 18528 34044 19552
rect 33724 18464 33732 18528
rect 33796 18464 33812 18528
rect 33876 18464 33892 18528
rect 33956 18464 33972 18528
rect 34036 18464 34044 18528
rect 33724 17440 34044 18464
rect 33724 17376 33732 17440
rect 33796 17376 33812 17440
rect 33876 17376 33892 17440
rect 33956 17376 33972 17440
rect 34036 17376 34044 17440
rect 33724 16352 34044 17376
rect 33724 16288 33732 16352
rect 33796 16288 33812 16352
rect 33876 16288 33892 16352
rect 33956 16288 33972 16352
rect 34036 16288 34044 16352
rect 33724 15264 34044 16288
rect 33724 15200 33732 15264
rect 33796 15200 33812 15264
rect 33876 15200 33892 15264
rect 33956 15200 33972 15264
rect 34036 15200 34044 15264
rect 33724 14176 34044 15200
rect 33724 14112 33732 14176
rect 33796 14112 33812 14176
rect 33876 14112 33892 14176
rect 33956 14112 33972 14176
rect 34036 14112 34044 14176
rect 33724 13088 34044 14112
rect 33724 13024 33732 13088
rect 33796 13024 33812 13088
rect 33876 13024 33892 13088
rect 33956 13024 33972 13088
rect 34036 13024 34044 13088
rect 33724 12000 34044 13024
rect 33724 11936 33732 12000
rect 33796 11936 33812 12000
rect 33876 11936 33892 12000
rect 33956 11936 33972 12000
rect 34036 11936 34044 12000
rect 33724 10912 34044 11936
rect 33724 10848 33732 10912
rect 33796 10848 33812 10912
rect 33876 10848 33892 10912
rect 33956 10848 33972 10912
rect 34036 10848 34044 10912
rect 33724 9824 34044 10848
rect 33724 9760 33732 9824
rect 33796 9760 33812 9824
rect 33876 9760 33892 9824
rect 33956 9760 33972 9824
rect 34036 9760 34044 9824
rect 33724 8736 34044 9760
rect 33724 8672 33732 8736
rect 33796 8672 33812 8736
rect 33876 8672 33892 8736
rect 33956 8672 33972 8736
rect 34036 8672 34044 8736
rect 33724 7648 34044 8672
rect 33724 7584 33732 7648
rect 33796 7584 33812 7648
rect 33876 7584 33892 7648
rect 33956 7584 33972 7648
rect 34036 7584 34044 7648
rect 33724 6560 34044 7584
rect 33724 6496 33732 6560
rect 33796 6496 33812 6560
rect 33876 6496 33892 6560
rect 33956 6496 33972 6560
rect 34036 6496 34044 6560
rect 33724 5472 34044 6496
rect 33724 5408 33732 5472
rect 33796 5408 33812 5472
rect 33876 5408 33892 5472
rect 33956 5408 33972 5472
rect 34036 5408 34044 5472
rect 33724 4384 34044 5408
rect 33724 4320 33732 4384
rect 33796 4354 33812 4384
rect 33876 4354 33892 4384
rect 33956 4354 33972 4384
rect 34036 4320 34044 4384
rect 33724 4118 33766 4320
rect 34002 4118 34044 4320
rect 33724 3296 34044 4118
rect 33724 3232 33732 3296
rect 33796 3232 33812 3296
rect 33876 3232 33892 3296
rect 33956 3232 33972 3296
rect 34036 3232 34044 3296
rect 33724 2208 34044 3232
rect 33724 2144 33732 2208
rect 33796 2144 33812 2208
rect 33876 2144 33892 2208
rect 33956 2144 33972 2208
rect 34036 2144 34044 2208
rect 33724 2128 34044 2144
<< via4 >>
rect 2386 34304 2622 34330
rect 2386 34240 2416 34304
rect 2416 34240 2432 34304
rect 2432 34240 2496 34304
rect 2496 34240 2512 34304
rect 2512 34240 2576 34304
rect 2576 34240 2592 34304
rect 2592 34240 2622 34304
rect 2386 34094 2622 34240
rect 2386 3458 2622 3694
rect 3046 34848 3282 34990
rect 3046 34784 3076 34848
rect 3076 34784 3092 34848
rect 3092 34784 3156 34848
rect 3156 34784 3172 34848
rect 3172 34784 3236 34848
rect 3236 34784 3252 34848
rect 3252 34784 3282 34848
rect 3046 34754 3282 34784
rect 3046 4320 3076 4354
rect 3076 4320 3092 4354
rect 3092 4320 3156 4354
rect 3156 4320 3172 4354
rect 3172 4320 3236 4354
rect 3236 4320 3252 4354
rect 3252 4320 3282 4354
rect 3046 4118 3282 4320
rect 33106 34304 33342 34330
rect 33106 34240 33136 34304
rect 33136 34240 33152 34304
rect 33152 34240 33216 34304
rect 33216 34240 33232 34304
rect 33232 34240 33296 34304
rect 33296 34240 33312 34304
rect 33312 34240 33342 34304
rect 33106 34094 33342 34240
rect 33106 3458 33342 3694
rect 33766 34848 34002 34990
rect 33766 34784 33796 34848
rect 33796 34784 33812 34848
rect 33812 34784 33876 34848
rect 33876 34784 33892 34848
rect 33892 34784 33956 34848
rect 33956 34784 33972 34848
rect 33972 34784 34002 34848
rect 33766 34754 34002 34784
rect 33766 4320 33796 4354
rect 33796 4320 33812 4354
rect 33812 4320 33876 4354
rect 33876 4320 33892 4354
rect 33892 4320 33956 4354
rect 33956 4320 33972 4354
rect 33972 4320 34002 4354
rect 33766 4118 34002 4320
<< metal5 >>
rect 1056 34990 58928 35032
rect 1056 34754 3046 34990
rect 3282 34754 33766 34990
rect 34002 34754 58928 34990
rect 1056 34712 58928 34754
rect 1056 34330 58928 34372
rect 1056 34094 2386 34330
rect 2622 34094 33106 34330
rect 33342 34094 58928 34330
rect 1056 34052 58928 34094
rect 1056 4354 58928 4396
rect 1056 4118 3046 4354
rect 3282 4118 33766 4354
rect 34002 4118 58928 4354
rect 1056 4076 58928 4118
rect 1056 3694 58928 3736
rect 1056 3458 2386 3694
rect 2622 3458 33106 3694
rect 33342 3458 58928 3694
rect 1056 3416 58928 3458
use sky130_fd_sc_hd__buf_4  _063_
timestamp 0
transform 1 0 17756 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _064_
timestamp 0
transform 1 0 32108 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp 0
transform -1 0 32016 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _066_
timestamp 0
transform -1 0 34776 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 0
transform 1 0 34776 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _068_
timestamp 0
transform -1 0 37168 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 0
transform -1 0 37536 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _070_
timestamp 0
transform -1 0 38916 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 0
transform 1 0 38916 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _072_
timestamp 0
transform 1 0 39836 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 0
transform -1 0 39836 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _074_
timestamp 0
transform 1 0 42412 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 0
transform -1 0 41768 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _076_
timestamp 0
transform 1 0 43240 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 0
transform 1 0 43240 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _078_
timestamp 0
transform -1 0 44896 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 0
transform -1 0 44620 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _080_
timestamp 0
transform 1 0 44896 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 0
transform 1 0 44620 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _082_
timestamp 0
transform -1 0 17204 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _083_
timestamp 0
transform -1 0 49772 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 0
transform 1 0 49772 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _085_
timestamp 0
transform -1 0 51888 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 0
transform 1 0 51888 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _087_
timestamp 0
transform -1 0 52532 0 1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 0
transform 1 0 52164 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _089_
timestamp 0
transform 1 0 52532 0 1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 0
transform -1 0 51060 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _091_
timestamp 0
transform 1 0 52716 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 0
transform -1 0 51704 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _093_
timestamp 0
transform -1 0 19688 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 0
transform -1 0 19136 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _095_
timestamp 0
transform 1 0 16560 0 1 55488
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 0
transform -1 0 16928 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _097_
timestamp 0
transform 1 0 16928 0 1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 0
transform -1 0 16560 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _099_
timestamp 0
transform 1 0 15824 0 1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 0
transform -1 0 15824 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _101_
timestamp 0
transform -1 0 15732 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 0
transform -1 0 16008 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _103_
timestamp 0
transform 1 0 15732 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 0
transform -1 0 16284 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _105_
timestamp 0
transform 1 0 16836 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _106_
timestamp 0
transform -1 0 18216 0 1 55488
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 0
transform -1 0 18584 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _108_
timestamp 0
transform 1 0 17388 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 0
transform -1 0 17756 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _110_
timestamp 0
transform 1 0 18216 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 0
transform -1 0 18584 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _112_
timestamp 0
transform -1 0 19872 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 0
transform -1 0 19964 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _114_
timestamp 0
transform -1 0 22632 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 0
transform 1 0 22632 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _116_
timestamp 0
transform -1 0 24012 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 0
transform 1 0 24012 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _118_
timestamp 0
transform -1 0 25668 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 0
transform 1 0 25668 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _120_
timestamp 0
transform -1 0 26864 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 0
transform 1 0 26956 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _122_
timestamp 0
transform -1 0 28244 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 0
transform 1 0 27968 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _124_
timestamp 0
transform 1 0 28244 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 0
transform -1 0 28336 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _126_
timestamp 0
transform 1 0 32108 0 -1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _127_
timestamp 0
transform 1 0 33948 0 -1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _128_
timestamp 0
transform -1 0 38088 0 1 54400
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _129_
timestamp 0
transform 1 0 37996 0 -1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _130_
timestamp 0
transform 1 0 39836 0 -1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _131_
timestamp 0
transform 1 0 41676 0 1 54400
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _132_
timestamp 0
transform 1 0 42964 0 -1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _133_
timestamp 0
transform 1 0 44804 0 -1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _134_
timestamp 0
transform 1 0 44068 0 -1 54400
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _135_
timestamp 0
transform 1 0 48852 0 -1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _136_
timestamp 0
transform 1 0 50784 0 -1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _137_
timestamp 0
transform 1 0 51336 0 1 54400
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _138_
timestamp 0
transform 1 0 52716 0 -1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _139_
timestamp 0
transform 1 0 51336 0 1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _140_
timestamp 0
transform -1 0 24748 0 -1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _141_
timestamp 0
transform -1 0 21712 0 -1 56576
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _142_
timestamp 0
transform -1 0 19872 0 -1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _143_
timestamp 0
transform -1 0 21712 0 -1 54400
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _144_
timestamp 0
transform -1 0 22448 0 1 54400
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _145_
timestamp 0
transform -1 0 22264 0 1 56576
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _146_
timestamp 0
transform -1 0 22540 0 1 53312
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _147_
timestamp 0
transform -1 0 21712 0 -1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _148_
timestamp 0
transform 1 0 22448 0 1 54400
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _149_
timestamp 0
transform -1 0 21436 0 -1 53312
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _150_
timestamp 0
transform 1 0 20608 0 1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _151_
timestamp 0
transform 1 0 22448 0 1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _152_
timestamp 0
transform 1 0 24748 0 -1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _153_
timestamp 0
transform 1 0 26220 0 1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _154_
timestamp 0
transform 1 0 27600 0 1 54400
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _155_
timestamp 0
transform 1 0 28152 0 -1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform -1 0 38088 0 1 55488
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 0
transform -1 0 27600 0 1 54400
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 0
transform -1 0 27876 0 1 53312
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 0
transform 1 0 39836 0 1 54400
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 0
transform 1 0 44988 0 1 54400
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout1
timestamp 0
transform -1 0 24932 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout2
timestamp 0
transform -1 0 35696 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout3
timestamp 0
transform -1 0 53728 0 1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 0
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 0
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 0
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 0
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 0
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 0
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 0
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 0
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 0
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 0
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 0
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 0
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 0
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 0
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 0
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 0
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 0
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 0
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 0
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 0
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 0
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 0
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 0
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 0
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 0
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 0
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 0
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 0
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_365
timestamp 0
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_377
timestamp 0
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 0
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_393
timestamp 0
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_405
timestamp 0
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_417
timestamp 0
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_421
timestamp 0
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_433
timestamp 0
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_445
timestamp 0
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_449
timestamp 0
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_461
timestamp 0
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_473
timestamp 0
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_477
timestamp 0
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_489
timestamp 0
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_501
timestamp 0
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_505
timestamp 0
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_517
timestamp 0
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_529
timestamp 0
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_533
timestamp 0
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_545
timestamp 0
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_557
timestamp 0
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_561
timestamp 0
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_573
timestamp 0
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_585
timestamp 0
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_589
timestamp 0
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_601
timestamp 0
transform 1 0 56396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_613
timestamp 0
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_617
timestamp 0
transform 1 0 57868 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 0
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 0
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 0
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 0
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 0
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 0
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 0
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 0
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 0
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 0
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 0
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 0
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 0
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 0
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 0
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 0
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 0
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 0
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 0
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 0
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 0
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 0
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 0
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 0
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 0
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 0
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 0
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 0
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 0
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 0
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 0
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 0
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 0
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 0
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_385
timestamp 0
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 0
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_393
timestamp 0
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_405
timestamp 0
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_417
timestamp 0
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_429
timestamp 0
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_441
timestamp 0
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_447
timestamp 0
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_449
timestamp 0
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_461
timestamp 0
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_473
timestamp 0
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_485
timestamp 0
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_497
timestamp 0
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_503
timestamp 0
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_505
timestamp 0
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_517
timestamp 0
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_529
timestamp 0
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_541
timestamp 0
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_553
timestamp 0
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_559
timestamp 0
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_561
timestamp 0
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_573
timestamp 0
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_585
timestamp 0
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_597
timestamp 0
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_609
timestamp 0
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_615
timestamp 0
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_617
timestamp 0
transform 1 0 57868 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 0
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 0
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 0
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 0
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 0
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 0
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 0
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 0
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 0
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 0
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 0
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 0
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 0
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 0
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 0
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 0
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 0
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 0
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 0
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 0
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 0
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 0
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 0
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 0
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 0
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 0
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 0
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 0
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 0
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 0
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 0
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 0
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 0
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 0
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 0
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 0
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_401
timestamp 0
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_413
timestamp 0
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 0
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 0
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 0
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_445
timestamp 0
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_457
timestamp 0
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_469
timestamp 0
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_475
timestamp 0
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_477
timestamp 0
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_489
timestamp 0
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_501
timestamp 0
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_513
timestamp 0
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_525
timestamp 0
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_531
timestamp 0
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_533
timestamp 0
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_545
timestamp 0
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_557
timestamp 0
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_569
timestamp 0
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_581
timestamp 0
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_587
timestamp 0
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_589
timestamp 0
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_601
timestamp 0
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_613
timestamp 0
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 0
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 0
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 0
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 0
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 0
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 0
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 0
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 0
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 0
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 0
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 0
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 0
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 0
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 0
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 0
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 0
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 0
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 0
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 0
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 0
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 0
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 0
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 0
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 0
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 0
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 0
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 0
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 0
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 0
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 0
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 0
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 0
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 0
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 0
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 0
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 0
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 0
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 0
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 0
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 0
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_429
timestamp 0
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_441
timestamp 0
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 0
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 0
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_461
timestamp 0
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_473
timestamp 0
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_485
timestamp 0
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_497
timestamp 0
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_503
timestamp 0
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_505
timestamp 0
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_517
timestamp 0
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_529
timestamp 0
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_541
timestamp 0
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_553
timestamp 0
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_559
timestamp 0
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_561
timestamp 0
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_573
timestamp 0
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_585
timestamp 0
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_597
timestamp 0
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_609
timestamp 0
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_615
timestamp 0
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_617
timestamp 0
transform 1 0 57868 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 0
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 0
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 0
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 0
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 0
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 0
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 0
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 0
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 0
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 0
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 0
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 0
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 0
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 0
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 0
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 0
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 0
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 0
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 0
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 0
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 0
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 0
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 0
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 0
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 0
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 0
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 0
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 0
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 0
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 0
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 0
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 0
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 0
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 0
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 0
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 0
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 0
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 0
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 0
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 0
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 0
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_457
timestamp 0
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_469
timestamp 0
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_475
timestamp 0
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_477
timestamp 0
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_489
timestamp 0
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_501
timestamp 0
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_513
timestamp 0
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_525
timestamp 0
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_531
timestamp 0
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_533
timestamp 0
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_545
timestamp 0
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_557
timestamp 0
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_569
timestamp 0
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_581
timestamp 0
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_587
timestamp 0
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_589
timestamp 0
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_601
timestamp 0
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_613
timestamp 0
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 0
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 0
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 0
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 0
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 0
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 0
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 0
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 0
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 0
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 0
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 0
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 0
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 0
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 0
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 0
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 0
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 0
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 0
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 0
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 0
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 0
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 0
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 0
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 0
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 0
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 0
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 0
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 0
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 0
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 0
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 0
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 0
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 0
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 0
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 0
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 0
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 0
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 0
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 0
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 0
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 0
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 0
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 0
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 0
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 0
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_461
timestamp 0
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_473
timestamp 0
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_485
timestamp 0
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_497
timestamp 0
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_503
timestamp 0
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_505
timestamp 0
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_517
timestamp 0
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_529
timestamp 0
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_541
timestamp 0
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_553
timestamp 0
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_559
timestamp 0
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_561
timestamp 0
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_573
timestamp 0
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_585
timestamp 0
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_597
timestamp 0
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_609
timestamp 0
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_615
timestamp 0
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_617
timestamp 0
transform 1 0 57868 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 0
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 0
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 0
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 0
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 0
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 0
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 0
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 0
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 0
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 0
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 0
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 0
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 0
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 0
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 0
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 0
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 0
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 0
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 0
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 0
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 0
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 0
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 0
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 0
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 0
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 0
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 0
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 0
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 0
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 0
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 0
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 0
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 0
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 0
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 0
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 0
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 0
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 0
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 0
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 0
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 0
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 0
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_457
timestamp 0
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_469
timestamp 0
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_475
timestamp 0
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_477
timestamp 0
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_489
timestamp 0
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_501
timestamp 0
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_513
timestamp 0
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_525
timestamp 0
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_531
timestamp 0
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_533
timestamp 0
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_545
timestamp 0
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_557
timestamp 0
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_569
timestamp 0
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_581
timestamp 0
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_587
timestamp 0
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_589
timestamp 0
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_601
timestamp 0
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_613
timestamp 0
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 0
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 0
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 0
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 0
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 0
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 0
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 0
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 0
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 0
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 0
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 0
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 0
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 0
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 0
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 0
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 0
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 0
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 0
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 0
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 0
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 0
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 0
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 0
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 0
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 0
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 0
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 0
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 0
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 0
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 0
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 0
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 0
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 0
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 0
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 0
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 0
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 0
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 0
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 0
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 0
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 0
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_429
timestamp 0
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_441
timestamp 0
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 0
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_449
timestamp 0
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_461
timestamp 0
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_473
timestamp 0
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_485
timestamp 0
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_497
timestamp 0
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_503
timestamp 0
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_505
timestamp 0
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_517
timestamp 0
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_529
timestamp 0
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_541
timestamp 0
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_553
timestamp 0
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_559
timestamp 0
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_561
timestamp 0
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_573
timestamp 0
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_585
timestamp 0
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_597
timestamp 0
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_609
timestamp 0
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_615
timestamp 0
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_617
timestamp 0
transform 1 0 57868 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 0
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 0
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 0
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 0
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 0
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 0
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 0
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 0
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 0
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 0
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 0
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 0
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 0
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 0
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 0
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 0
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 0
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 0
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 0
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 0
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 0
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 0
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 0
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 0
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 0
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 0
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 0
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 0
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 0
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 0
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 0
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 0
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 0
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 0
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 0
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_401
timestamp 0
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_413
timestamp 0
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 0
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 0
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 0
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 0
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_457
timestamp 0
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_469
timestamp 0
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_475
timestamp 0
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_477
timestamp 0
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_489
timestamp 0
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_501
timestamp 0
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_513
timestamp 0
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_525
timestamp 0
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_531
timestamp 0
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_533
timestamp 0
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_545
timestamp 0
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_557
timestamp 0
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_569
timestamp 0
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_581
timestamp 0
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_587
timestamp 0
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_589
timestamp 0
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_601
timestamp 0
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_613
timestamp 0
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 0
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 0
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 0
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 0
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 0
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 0
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 0
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 0
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 0
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 0
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 0
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 0
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 0
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 0
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 0
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 0
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 0
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 0
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 0
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 0
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 0
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 0
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 0
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 0
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 0
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 0
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 0
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 0
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 0
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 0
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 0
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 0
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 0
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 0
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 0
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 0
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 0
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 0
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 0
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 0
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_405
timestamp 0
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_417
timestamp 0
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_429
timestamp 0
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_441
timestamp 0
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_447
timestamp 0
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_449
timestamp 0
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_461
timestamp 0
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_473
timestamp 0
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_485
timestamp 0
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_497
timestamp 0
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_503
timestamp 0
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_505
timestamp 0
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_517
timestamp 0
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_529
timestamp 0
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_541
timestamp 0
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_553
timestamp 0
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_559
timestamp 0
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_561
timestamp 0
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_573
timestamp 0
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_585
timestamp 0
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_597
timestamp 0
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_609
timestamp 0
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_615
timestamp 0
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_617
timestamp 0
transform 1 0 57868 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 0
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 0
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 0
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 0
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 0
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 0
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 0
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 0
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 0
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 0
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 0
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 0
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 0
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 0
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 0
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 0
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 0
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 0
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 0
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 0
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 0
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 0
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 0
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 0
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 0
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 0
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 0
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 0
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 0
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 0
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 0
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 0
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 0
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 0
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 0
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 0
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 0
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 0
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 0
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_401
timestamp 0
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_413
timestamp 0
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_419
timestamp 0
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_421
timestamp 0
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_433
timestamp 0
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_445
timestamp 0
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_457
timestamp 0
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_469
timestamp 0
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_475
timestamp 0
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_477
timestamp 0
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_489
timestamp 0
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_501
timestamp 0
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_513
timestamp 0
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_525
timestamp 0
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_531
timestamp 0
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_533
timestamp 0
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_545
timestamp 0
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_557
timestamp 0
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_569
timestamp 0
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_581
timestamp 0
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_587
timestamp 0
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_589
timestamp 0
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_601
timestamp 0
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_613
timestamp 0
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 0
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 0
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 0
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 0
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 0
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 0
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 0
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 0
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 0
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 0
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 0
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 0
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 0
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 0
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 0
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 0
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 0
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 0
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 0
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 0
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 0
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 0
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 0
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 0
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 0
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 0
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 0
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 0
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 0
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 0
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 0
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 0
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 0
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 0
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 0
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 0
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 0
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 0
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 0
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_405
timestamp 0
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_417
timestamp 0
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_429
timestamp 0
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_441
timestamp 0
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 0
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_449
timestamp 0
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_461
timestamp 0
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_473
timestamp 0
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_485
timestamp 0
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_497
timestamp 0
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_503
timestamp 0
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_505
timestamp 0
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_517
timestamp 0
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_529
timestamp 0
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_541
timestamp 0
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_553
timestamp 0
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_559
timestamp 0
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_561
timestamp 0
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_573
timestamp 0
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_585
timestamp 0
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_597
timestamp 0
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_609
timestamp 0
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_615
timestamp 0
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_617
timestamp 0
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 0
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 0
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 0
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 0
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 0
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 0
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 0
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 0
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 0
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 0
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 0
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 0
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 0
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 0
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 0
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 0
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 0
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 0
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 0
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 0
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 0
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 0
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 0
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 0
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 0
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 0
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 0
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 0
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 0
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 0
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 0
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 0
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 0
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 0
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 0
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 0
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 0
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_389
timestamp 0
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_401
timestamp 0
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_413
timestamp 0
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_419
timestamp 0
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_421
timestamp 0
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_433
timestamp 0
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_445
timestamp 0
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_457
timestamp 0
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_469
timestamp 0
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_475
timestamp 0
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_477
timestamp 0
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_489
timestamp 0
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_501
timestamp 0
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_513
timestamp 0
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_525
timestamp 0
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_531
timestamp 0
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_533
timestamp 0
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_545
timestamp 0
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_557
timestamp 0
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_569
timestamp 0
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_581
timestamp 0
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_587
timestamp 0
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_589
timestamp 0
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_601
timestamp 0
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_613
timestamp 0
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 0
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 0
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 0
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 0
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 0
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 0
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 0
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 0
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 0
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 0
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 0
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 0
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 0
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 0
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 0
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 0
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 0
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 0
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 0
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 0
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 0
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 0
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 0
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 0
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 0
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 0
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 0
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 0
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 0
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 0
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 0
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_329
timestamp 0
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 0
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_337
timestamp 0
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_349
timestamp 0
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_361
timestamp 0
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_373
timestamp 0
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_385
timestamp 0
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_391
timestamp 0
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_393
timestamp 0
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_405
timestamp 0
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_417
timestamp 0
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_429
timestamp 0
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_441
timestamp 0
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_447
timestamp 0
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_449
timestamp 0
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_461
timestamp 0
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_473
timestamp 0
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_485
timestamp 0
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_497
timestamp 0
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_503
timestamp 0
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_505
timestamp 0
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_517
timestamp 0
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_529
timestamp 0
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_541
timestamp 0
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_553
timestamp 0
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_559
timestamp 0
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_561
timestamp 0
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_573
timestamp 0
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_585
timestamp 0
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_597
timestamp 0
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_609
timestamp 0
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_615
timestamp 0
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_617
timestamp 0
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 0
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 0
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 0
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 0
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 0
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 0
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 0
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 0
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 0
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 0
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 0
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 0
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 0
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 0
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 0
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 0
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 0
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 0
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 0
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 0
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_233
timestamp 0
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_245
timestamp 0
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 0
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 0
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 0
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 0
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_289
timestamp 0
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_301
timestamp 0
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 0
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 0
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_321
timestamp 0
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_333
timestamp 0
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_345
timestamp 0
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_357
timestamp 0
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_363
timestamp 0
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_365
timestamp 0
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_377
timestamp 0
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_389
timestamp 0
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_401
timestamp 0
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_413
timestamp 0
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_419
timestamp 0
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_421
timestamp 0
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_433
timestamp 0
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_445
timestamp 0
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_457
timestamp 0
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_469
timestamp 0
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_475
timestamp 0
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_477
timestamp 0
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_489
timestamp 0
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_501
timestamp 0
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_513
timestamp 0
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_525
timestamp 0
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_531
timestamp 0
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_533
timestamp 0
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_545
timestamp 0
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_557
timestamp 0
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_569
timestamp 0
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_581
timestamp 0
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_587
timestamp 0
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_589
timestamp 0
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_601
timestamp 0
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_613
timestamp 0
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 0
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 0
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 0
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 0
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 0
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 0
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 0
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 0
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 0
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 0
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 0
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 0
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 0
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 0
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 0
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 0
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 0
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_193
timestamp 0
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 0
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_217
timestamp 0
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 0
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 0
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 0
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_249
timestamp 0
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_261
timestamp 0
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_273
timestamp 0
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 0
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 0
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 0
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 0
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_317
timestamp 0
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_329
timestamp 0
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_335
timestamp 0
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_337
timestamp 0
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_349
timestamp 0
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_361
timestamp 0
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_373
timestamp 0
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_385
timestamp 0
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_391
timestamp 0
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_393
timestamp 0
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_405
timestamp 0
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_417
timestamp 0
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_429
timestamp 0
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_441
timestamp 0
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_447
timestamp 0
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_449
timestamp 0
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_461
timestamp 0
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_473
timestamp 0
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_485
timestamp 0
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_497
timestamp 0
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_503
timestamp 0
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_505
timestamp 0
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_517
timestamp 0
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_529
timestamp 0
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_541
timestamp 0
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_553
timestamp 0
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_559
timestamp 0
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_561
timestamp 0
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_573
timestamp 0
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_585
timestamp 0
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_597
timestamp 0
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_609
timestamp 0
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_615
timestamp 0
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_617
timestamp 0
transform 1 0 57868 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 0
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 0
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 0
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 0
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 0
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 0
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 0
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 0
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 0
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 0
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 0
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 0
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 0
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 0
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 0
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 0
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 0
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 0
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 0
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 0
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_221
timestamp 0
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_233
timestamp 0
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_245
timestamp 0
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 0
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 0
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 0
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 0
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 0
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 0
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 0
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 0
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_321
timestamp 0
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_333
timestamp 0
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_345
timestamp 0
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_357
timestamp 0
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_363
timestamp 0
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_365
timestamp 0
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_377
timestamp 0
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_389
timestamp 0
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_401
timestamp 0
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_413
timestamp 0
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_419
timestamp 0
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_421
timestamp 0
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_433
timestamp 0
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_445
timestamp 0
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_457
timestamp 0
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_469
timestamp 0
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_475
timestamp 0
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_477
timestamp 0
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_489
timestamp 0
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_501
timestamp 0
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_513
timestamp 0
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_525
timestamp 0
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_531
timestamp 0
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_533
timestamp 0
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_545
timestamp 0
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_557
timestamp 0
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_569
timestamp 0
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_581
timestamp 0
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_587
timestamp 0
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_589
timestamp 0
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_601
timestamp 0
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_613
timestamp 0
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 0
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 0
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 0
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 0
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 0
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 0
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 0
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 0
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 0
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 0
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 0
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 0
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 0
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 0
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 0
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 0
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 0
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_193
timestamp 0
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_205
timestamp 0
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 0
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 0
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 0
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 0
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 0
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 0
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 0
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 0
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 0
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 0
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 0
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 0
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_329
timestamp 0
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_335
timestamp 0
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_337
timestamp 0
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_349
timestamp 0
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_361
timestamp 0
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_373
timestamp 0
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_385
timestamp 0
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_391
timestamp 0
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_393
timestamp 0
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_405
timestamp 0
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_417
timestamp 0
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_429
timestamp 0
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_441
timestamp 0
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_447
timestamp 0
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_449
timestamp 0
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_461
timestamp 0
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_473
timestamp 0
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_485
timestamp 0
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_497
timestamp 0
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_503
timestamp 0
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_505
timestamp 0
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_517
timestamp 0
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_529
timestamp 0
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_541
timestamp 0
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_553
timestamp 0
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_559
timestamp 0
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_561
timestamp 0
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_573
timestamp 0
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_585
timestamp 0
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_597
timestamp 0
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_609
timestamp 0
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_615
timestamp 0
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_617
timestamp 0
transform 1 0 57868 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 0
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 0
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 0
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 0
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 0
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 0
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 0
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 0
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 0
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 0
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 0
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 0
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 0
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_165
timestamp 0
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 0
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_189
timestamp 0
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 0
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 0
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_209
timestamp 0
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_221
timestamp 0
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_233
timestamp 0
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_245
timestamp 0
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 0
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 0
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 0
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 0
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 0
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_301
timestamp 0
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 0
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 0
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_321
timestamp 0
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_333
timestamp 0
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_345
timestamp 0
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_357
timestamp 0
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_363
timestamp 0
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_365
timestamp 0
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_377
timestamp 0
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_389
timestamp 0
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_401
timestamp 0
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_413
timestamp 0
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_419
timestamp 0
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_421
timestamp 0
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_433
timestamp 0
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_445
timestamp 0
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_457
timestamp 0
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_469
timestamp 0
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_475
timestamp 0
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_477
timestamp 0
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_489
timestamp 0
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_501
timestamp 0
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_513
timestamp 0
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_525
timestamp 0
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_531
timestamp 0
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_533
timestamp 0
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_545
timestamp 0
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_557
timestamp 0
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_569
timestamp 0
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_581
timestamp 0
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_587
timestamp 0
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_589
timestamp 0
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_601
timestamp 0
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_613
timestamp 0
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 0
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 0
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 0
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 0
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 0
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 0
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 0
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 0
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 0
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 0
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 0
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 0
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 0
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 0
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 0
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 0
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 0
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_193
timestamp 0
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_205
timestamp 0
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_217
timestamp 0
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 0
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 0
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_237
timestamp 0
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_249
timestamp 0
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_261
timestamp 0
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_273
timestamp 0
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 0
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 0
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 0
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 0
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_317
timestamp 0
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_329
timestamp 0
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_335
timestamp 0
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_337
timestamp 0
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_349
timestamp 0
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_361
timestamp 0
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_373
timestamp 0
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_385
timestamp 0
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_391
timestamp 0
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_393
timestamp 0
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_405
timestamp 0
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_417
timestamp 0
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_429
timestamp 0
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_441
timestamp 0
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_447
timestamp 0
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_449
timestamp 0
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_461
timestamp 0
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_473
timestamp 0
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_485
timestamp 0
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_497
timestamp 0
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_503
timestamp 0
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_505
timestamp 0
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_517
timestamp 0
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_529
timestamp 0
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_541
timestamp 0
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_553
timestamp 0
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_559
timestamp 0
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_561
timestamp 0
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_573
timestamp 0
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_585
timestamp 0
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_597
timestamp 0
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_609
timestamp 0
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_615
timestamp 0
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_617
timestamp 0
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 0
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 0
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 0
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 0
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 0
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 0
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 0
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 0
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 0
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 0
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 0
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 0
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 0
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 0
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 0
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 0
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 0
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 0
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 0
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 0
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_221
timestamp 0
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_233
timestamp 0
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_245
timestamp 0
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 0
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 0
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 0
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_277
timestamp 0
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_289
timestamp 0
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_301
timestamp 0
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 0
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 0
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_321
timestamp 0
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_333
timestamp 0
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_345
timestamp 0
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_357
timestamp 0
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_363
timestamp 0
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_365
timestamp 0
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_377
timestamp 0
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_389
timestamp 0
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_401
timestamp 0
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_413
timestamp 0
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_419
timestamp 0
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_421
timestamp 0
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_433
timestamp 0
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_445
timestamp 0
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_457
timestamp 0
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_469
timestamp 0
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_475
timestamp 0
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_477
timestamp 0
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_489
timestamp 0
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_501
timestamp 0
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_513
timestamp 0
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_525
timestamp 0
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_531
timestamp 0
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_533
timestamp 0
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_545
timestamp 0
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_557
timestamp 0
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_569
timestamp 0
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_581
timestamp 0
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_587
timestamp 0
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_589
timestamp 0
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_601
timestamp 0
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_613
timestamp 0
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 0
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 0
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 0
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 0
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 0
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 0
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 0
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 0
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 0
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 0
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 0
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 0
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 0
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 0
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 0
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 0
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 0
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 0
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_193
timestamp 0
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_205
timestamp 0
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_217
timestamp 0
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 0
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 0
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 0
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 0
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 0
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_273
timestamp 0
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 0
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 0
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 0
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 0
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_317
timestamp 0
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_329
timestamp 0
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_335
timestamp 0
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_337
timestamp 0
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_349
timestamp 0
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_361
timestamp 0
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_373
timestamp 0
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_385
timestamp 0
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_391
timestamp 0
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_393
timestamp 0
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_405
timestamp 0
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_417
timestamp 0
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_429
timestamp 0
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_441
timestamp 0
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_447
timestamp 0
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_449
timestamp 0
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_461
timestamp 0
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_473
timestamp 0
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_485
timestamp 0
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_497
timestamp 0
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_503
timestamp 0
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_505
timestamp 0
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_517
timestamp 0
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_529
timestamp 0
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_541
timestamp 0
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_553
timestamp 0
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_559
timestamp 0
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_561
timestamp 0
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_573
timestamp 0
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_585
timestamp 0
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_597
timestamp 0
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_609
timestamp 0
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_615
timestamp 0
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_617
timestamp 0
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 0
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 0
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 0
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 0
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 0
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 0
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 0
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 0
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 0
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 0
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 0
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 0
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 0
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 0
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 0
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 0
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 0
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 0
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 0
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 0
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_221
timestamp 0
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_233
timestamp 0
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_245
timestamp 0
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 0
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 0
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 0
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 0
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 0
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 0
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 0
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 0
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_321
timestamp 0
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_333
timestamp 0
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_345
timestamp 0
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_357
timestamp 0
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_363
timestamp 0
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_365
timestamp 0
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_377
timestamp 0
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_389
timestamp 0
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_401
timestamp 0
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_413
timestamp 0
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_419
timestamp 0
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_421
timestamp 0
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_433
timestamp 0
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_445
timestamp 0
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_457
timestamp 0
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_469
timestamp 0
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_475
timestamp 0
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_477
timestamp 0
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_489
timestamp 0
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_501
timestamp 0
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_513
timestamp 0
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_525
timestamp 0
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_531
timestamp 0
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_533
timestamp 0
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_545
timestamp 0
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_557
timestamp 0
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_569
timestamp 0
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_581
timestamp 0
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_587
timestamp 0
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_589
timestamp 0
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_601
timestamp 0
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_613
timestamp 0
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 0
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 0
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 0
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 0
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 0
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 0
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 0
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 0
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 0
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 0
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 0
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 0
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 0
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 0
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 0
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 0
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 0
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 0
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_193
timestamp 0
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_205
timestamp 0
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 0
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 0
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 0
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 0
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 0
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_261
timestamp 0
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp 0
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 0
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 0
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 0
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 0
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_317
timestamp 0
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_329
timestamp 0
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_335
timestamp 0
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_337
timestamp 0
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_349
timestamp 0
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_361
timestamp 0
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_373
timestamp 0
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_385
timestamp 0
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_391
timestamp 0
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_393
timestamp 0
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_405
timestamp 0
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_417
timestamp 0
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_429
timestamp 0
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_441
timestamp 0
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_447
timestamp 0
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_449
timestamp 0
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_461
timestamp 0
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_473
timestamp 0
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_485
timestamp 0
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_497
timestamp 0
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_503
timestamp 0
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_505
timestamp 0
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_517
timestamp 0
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_529
timestamp 0
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_541
timestamp 0
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_553
timestamp 0
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_559
timestamp 0
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_561
timestamp 0
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_573
timestamp 0
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_585
timestamp 0
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_597
timestamp 0
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_609
timestamp 0
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_615
timestamp 0
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_617
timestamp 0
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 0
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 0
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 0
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 0
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 0
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 0
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 0
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 0
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 0
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 0
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 0
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 0
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 0
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 0
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 0
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 0
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 0
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 0
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 0
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 0
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 0
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_209
timestamp 0
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_221
timestamp 0
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_233
timestamp 0
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp 0
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 0
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 0
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 0
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_277
timestamp 0
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_289
timestamp 0
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 0
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 0
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 0
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_321
timestamp 0
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_333
timestamp 0
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_345
timestamp 0
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_357
timestamp 0
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_363
timestamp 0
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_365
timestamp 0
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_377
timestamp 0
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_389
timestamp 0
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_401
timestamp 0
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_413
timestamp 0
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_419
timestamp 0
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_421
timestamp 0
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_433
timestamp 0
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_445
timestamp 0
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_457
timestamp 0
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_469
timestamp 0
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_475
timestamp 0
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_477
timestamp 0
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_489
timestamp 0
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_501
timestamp 0
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_513
timestamp 0
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_525
timestamp 0
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_531
timestamp 0
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_533
timestamp 0
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_545
timestamp 0
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_557
timestamp 0
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_569
timestamp 0
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_581
timestamp 0
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_587
timestamp 0
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_589
timestamp 0
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_601
timestamp 0
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_613
timestamp 0
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 0
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 0
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 0
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 0
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 0
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 0
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 0
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 0
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 0
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 0
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 0
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 0
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 0
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 0
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 0
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 0
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 0
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 0
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 0
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 0
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 0
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 0
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 0
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 0
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 0
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 0
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_249
timestamp 0
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_261
timestamp 0
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_273
timestamp 0
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 0
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 0
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 0
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 0
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_317
timestamp 0
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_329
timestamp 0
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_335
timestamp 0
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_337
timestamp 0
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_349
timestamp 0
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_361
timestamp 0
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_373
timestamp 0
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_385
timestamp 0
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_391
timestamp 0
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_393
timestamp 0
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_405
timestamp 0
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_417
timestamp 0
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_429
timestamp 0
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_441
timestamp 0
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_447
timestamp 0
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_449
timestamp 0
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_461
timestamp 0
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_473
timestamp 0
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_485
timestamp 0
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_497
timestamp 0
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_503
timestamp 0
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_505
timestamp 0
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_517
timestamp 0
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_529
timestamp 0
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_541
timestamp 0
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_553
timestamp 0
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_559
timestamp 0
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_561
timestamp 0
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_573
timestamp 0
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_585
timestamp 0
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_597
timestamp 0
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_609
timestamp 0
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_615
timestamp 0
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_617
timestamp 0
transform 1 0 57868 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 0
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 0
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 0
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 0
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 0
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 0
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 0
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 0
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 0
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 0
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 0
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 0
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 0
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 0
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 0
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 0
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 0
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 0
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 0
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 0
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 0
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 0
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 0
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 0
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_233
timestamp 0
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_245
timestamp 0
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 0
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 0
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 0
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 0
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 0
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 0
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 0
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 0
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_321
timestamp 0
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_333
timestamp 0
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_345
timestamp 0
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_357
timestamp 0
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_363
timestamp 0
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_365
timestamp 0
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_377
timestamp 0
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_389
timestamp 0
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_401
timestamp 0
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_413
timestamp 0
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_419
timestamp 0
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_421
timestamp 0
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_433
timestamp 0
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_445
timestamp 0
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_457
timestamp 0
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_469
timestamp 0
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_475
timestamp 0
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_477
timestamp 0
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_489
timestamp 0
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_501
timestamp 0
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_513
timestamp 0
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_525
timestamp 0
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_531
timestamp 0
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_533
timestamp 0
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_545
timestamp 0
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_557
timestamp 0
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_569
timestamp 0
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_581
timestamp 0
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_587
timestamp 0
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_589
timestamp 0
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_601
timestamp 0
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_613
timestamp 0
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 0
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 0
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 0
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 0
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 0
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 0
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 0
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 0
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 0
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 0
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 0
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 0
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 0
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 0
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 0
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 0
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 0
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 0
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 0
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 0
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_193
timestamp 0
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_205
timestamp 0
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 0
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 0
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 0
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 0
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 0
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_261
timestamp 0
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 0
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 0
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 0
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 0
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 0
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_317
timestamp 0
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_329
timestamp 0
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_335
timestamp 0
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_337
timestamp 0
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_349
timestamp 0
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_361
timestamp 0
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_373
timestamp 0
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_385
timestamp 0
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_391
timestamp 0
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_393
timestamp 0
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_405
timestamp 0
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_417
timestamp 0
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_429
timestamp 0
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_441
timestamp 0
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_447
timestamp 0
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_449
timestamp 0
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_461
timestamp 0
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_473
timestamp 0
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_485
timestamp 0
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_497
timestamp 0
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_503
timestamp 0
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_505
timestamp 0
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_517
timestamp 0
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_529
timestamp 0
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_541
timestamp 0
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_553
timestamp 0
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_559
timestamp 0
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_561
timestamp 0
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_573
timestamp 0
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_585
timestamp 0
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_597
timestamp 0
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_609
timestamp 0
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_615
timestamp 0
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_617
timestamp 0
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 0
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 0
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 0
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 0
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 0
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 0
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 0
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 0
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 0
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 0
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 0
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 0
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 0
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 0
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 0
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 0
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 0
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 0
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 0
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 0
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 0
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 0
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 0
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 0
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_233
timestamp 0
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 0
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 0
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 0
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 0
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 0
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_289
timestamp 0
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_301
timestamp 0
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 0
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 0
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_321
timestamp 0
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_333
timestamp 0
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_345
timestamp 0
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_357
timestamp 0
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_363
timestamp 0
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_365
timestamp 0
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_377
timestamp 0
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_389
timestamp 0
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_401
timestamp 0
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_413
timestamp 0
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_419
timestamp 0
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_421
timestamp 0
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_433
timestamp 0
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_445
timestamp 0
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_457
timestamp 0
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_469
timestamp 0
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_475
timestamp 0
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_477
timestamp 0
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_489
timestamp 0
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_501
timestamp 0
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_513
timestamp 0
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_525
timestamp 0
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_531
timestamp 0
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_533
timestamp 0
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_545
timestamp 0
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_557
timestamp 0
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_569
timestamp 0
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_581
timestamp 0
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_587
timestamp 0
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_589
timestamp 0
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_601
timestamp 0
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_613
timestamp 0
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 0
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 0
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 0
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 0
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 0
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 0
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 0
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 0
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 0
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 0
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 0
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 0
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 0
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 0
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 0
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 0
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 0
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 0
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 0
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 0
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_193
timestamp 0
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 0
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 0
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 0
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 0
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 0
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 0
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 0
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 0
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 0
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 0
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 0
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 0
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_317
timestamp 0
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_329
timestamp 0
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 0
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_337
timestamp 0
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_349
timestamp 0
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_361
timestamp 0
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_373
timestamp 0
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_385
timestamp 0
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_391
timestamp 0
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_393
timestamp 0
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_405
timestamp 0
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_417
timestamp 0
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_429
timestamp 0
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_441
timestamp 0
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_447
timestamp 0
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_449
timestamp 0
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_461
timestamp 0
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_473
timestamp 0
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_485
timestamp 0
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_497
timestamp 0
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_503
timestamp 0
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_505
timestamp 0
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_517
timestamp 0
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_529
timestamp 0
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_541
timestamp 0
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_553
timestamp 0
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_559
timestamp 0
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_561
timestamp 0
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_573
timestamp 0
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_585
timestamp 0
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_597
timestamp 0
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_609
timestamp 0
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_615
timestamp 0
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_617
timestamp 0
transform 1 0 57868 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 0
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 0
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 0
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 0
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 0
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 0
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 0
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 0
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 0
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 0
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 0
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 0
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 0
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 0
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 0
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 0
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 0
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 0
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 0
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 0
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 0
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 0
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 0
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 0
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 0
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 0
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 0
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 0
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 0
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 0
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 0
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_301
timestamp 0
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 0
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 0
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_321
timestamp 0
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_333
timestamp 0
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_345
timestamp 0
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_357
timestamp 0
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_363
timestamp 0
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_365
timestamp 0
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_377
timestamp 0
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_389
timestamp 0
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_401
timestamp 0
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_413
timestamp 0
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_419
timestamp 0
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_421
timestamp 0
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_433
timestamp 0
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_445
timestamp 0
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_457
timestamp 0
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_469
timestamp 0
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_475
timestamp 0
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_477
timestamp 0
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_489
timestamp 0
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_501
timestamp 0
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_513
timestamp 0
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_525
timestamp 0
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_531
timestamp 0
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_533
timestamp 0
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_545
timestamp 0
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_557
timestamp 0
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_569
timestamp 0
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_581
timestamp 0
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_587
timestamp 0
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_589
timestamp 0
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_601
timestamp 0
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_613
timestamp 0
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 0
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 0
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 0
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 0
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 0
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 0
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 0
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 0
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 0
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 0
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 0
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 0
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 0
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 0
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 0
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 0
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 0
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 0
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 0
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 0
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_193
timestamp 0
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_205
timestamp 0
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 0
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 0
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 0
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 0
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 0
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 0
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 0
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 0
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 0
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 0
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_305
timestamp 0
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 0
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_329
timestamp 0
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_335
timestamp 0
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_337
timestamp 0
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_349
timestamp 0
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_361
timestamp 0
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_373
timestamp 0
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_385
timestamp 0
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_391
timestamp 0
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_393
timestamp 0
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_405
timestamp 0
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_417
timestamp 0
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_429
timestamp 0
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_441
timestamp 0
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_447
timestamp 0
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_449
timestamp 0
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_461
timestamp 0
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_473
timestamp 0
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_485
timestamp 0
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_497
timestamp 0
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_503
timestamp 0
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_505
timestamp 0
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_517
timestamp 0
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_529
timestamp 0
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_541
timestamp 0
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_553
timestamp 0
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_559
timestamp 0
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_561
timestamp 0
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_573
timestamp 0
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_585
timestamp 0
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_597
timestamp 0
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_609
timestamp 0
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_615
timestamp 0
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_617
timestamp 0
transform 1 0 57868 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 0
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 0
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 0
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 0
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 0
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 0
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 0
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 0
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 0
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 0
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 0
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 0
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 0
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 0
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 0
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 0
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 0
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 0
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 0
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 0
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 0
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 0
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 0
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 0
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 0
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 0
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 0
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 0
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 0
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_277
timestamp 0
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_289
timestamp 0
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_301
timestamp 0
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 0
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 0
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_321
timestamp 0
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_333
timestamp 0
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_345
timestamp 0
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_357
timestamp 0
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_363
timestamp 0
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_365
timestamp 0
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_377
timestamp 0
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_389
timestamp 0
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_401
timestamp 0
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_413
timestamp 0
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_419
timestamp 0
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_421
timestamp 0
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_433
timestamp 0
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_445
timestamp 0
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_457
timestamp 0
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_469
timestamp 0
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_475
timestamp 0
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_477
timestamp 0
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_489
timestamp 0
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_501
timestamp 0
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_513
timestamp 0
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_525
timestamp 0
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_531
timestamp 0
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_533
timestamp 0
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_545
timestamp 0
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_557
timestamp 0
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_569
timestamp 0
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_581
timestamp 0
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_587
timestamp 0
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_589
timestamp 0
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_601
timestamp 0
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_613
timestamp 0
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 0
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 0
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 0
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 0
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 0
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 0
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 0
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 0
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 0
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 0
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_105
timestamp 0
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 0
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 0
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 0
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_137
timestamp 0
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_149
timestamp 0
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_161
timestamp 0
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 0
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 0
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 0
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_193
timestamp 0
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_205
timestamp 0
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_217
timestamp 0
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 0
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 0
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 0
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_249
timestamp 0
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_261
timestamp 0
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_273
timestamp 0
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 0
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 0
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 0
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_305
timestamp 0
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_317
timestamp 0
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_329
timestamp 0
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_335
timestamp 0
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_337
timestamp 0
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_349
timestamp 0
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_361
timestamp 0
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_373
timestamp 0
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_385
timestamp 0
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_391
timestamp 0
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_393
timestamp 0
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_405
timestamp 0
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_417
timestamp 0
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_429
timestamp 0
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_441
timestamp 0
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_447
timestamp 0
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_449
timestamp 0
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_461
timestamp 0
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_473
timestamp 0
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_485
timestamp 0
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_497
timestamp 0
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_503
timestamp 0
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_505
timestamp 0
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_517
timestamp 0
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_529
timestamp 0
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_541
timestamp 0
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_553
timestamp 0
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_559
timestamp 0
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_561
timestamp 0
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_573
timestamp 0
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_585
timestamp 0
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_597
timestamp 0
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_609
timestamp 0
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_615
timestamp 0
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_617
timestamp 0
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 0
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 0
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 0
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 0
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 0
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 0
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 0
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_77
timestamp 0
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 0
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 0
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_97
timestamp 0
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_109
timestamp 0
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_121
timestamp 0
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_133
timestamp 0
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 0
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 0
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_153
timestamp 0
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_165
timestamp 0
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_177
timestamp 0
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_189
timestamp 0
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 0
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 0
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_209
timestamp 0
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_221
timestamp 0
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_233
timestamp 0
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_245
timestamp 0
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 0
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 0
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_265
timestamp 0
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_277
timestamp 0
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_289
timestamp 0
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_301
timestamp 0
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_307
timestamp 0
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_309
timestamp 0
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_321
timestamp 0
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_333
timestamp 0
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_345
timestamp 0
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_357
timestamp 0
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_363
timestamp 0
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_365
timestamp 0
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_377
timestamp 0
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_389
timestamp 0
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_401
timestamp 0
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_413
timestamp 0
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_419
timestamp 0
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_421
timestamp 0
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_433
timestamp 0
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_445
timestamp 0
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_457
timestamp 0
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_469
timestamp 0
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_475
timestamp 0
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_477
timestamp 0
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_489
timestamp 0
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_501
timestamp 0
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_513
timestamp 0
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_525
timestamp 0
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_531
timestamp 0
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_533
timestamp 0
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_545
timestamp 0
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_557
timestamp 0
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_569
timestamp 0
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_581
timestamp 0
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_587
timestamp 0
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_589
timestamp 0
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_601
timestamp 0
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_613
timestamp 0
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 0
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 0
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 0
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 0
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 0
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 0
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 0
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 0
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_81
timestamp 0
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_93
timestamp 0
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_105
timestamp 0
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 0
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 0
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 0
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_137
timestamp 0
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_149
timestamp 0
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_161
timestamp 0
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 0
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 0
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_181
timestamp 0
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_193
timestamp 0
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_205
timestamp 0
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_217
timestamp 0
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 0
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 0
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_237
timestamp 0
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_249
timestamp 0
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_261
timestamp 0
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_273
timestamp 0
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 0
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 0
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_293
timestamp 0
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_305
timestamp 0
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_317
timestamp 0
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_329
timestamp 0
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_335
timestamp 0
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_337
timestamp 0
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_349
timestamp 0
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_361
timestamp 0
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_373
timestamp 0
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_385
timestamp 0
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_391
timestamp 0
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_393
timestamp 0
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_405
timestamp 0
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_417
timestamp 0
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_429
timestamp 0
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_441
timestamp 0
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_447
timestamp 0
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_449
timestamp 0
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_461
timestamp 0
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_473
timestamp 0
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_485
timestamp 0
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_497
timestamp 0
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_503
timestamp 0
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_505
timestamp 0
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_517
timestamp 0
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_529
timestamp 0
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_541
timestamp 0
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_553
timestamp 0
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_559
timestamp 0
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_561
timestamp 0
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_573
timestamp 0
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_585
timestamp 0
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_597
timestamp 0
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_609
timestamp 0
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_615
timestamp 0
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_617
timestamp 0
transform 1 0 57868 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 0
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 0
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 0
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 0
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 0
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 0
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 0
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 0
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 0
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 0
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 0
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 0
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 0
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 0
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 0
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 0
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_153
timestamp 0
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_165
timestamp 0
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_177
timestamp 0
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_189
timestamp 0
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 0
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 0
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_209
timestamp 0
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_221
timestamp 0
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_233
timestamp 0
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_245
timestamp 0
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 0
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 0
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_265
timestamp 0
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_277
timestamp 0
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_289
timestamp 0
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_301
timestamp 0
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 0
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 0
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_321
timestamp 0
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_333
timestamp 0
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_345
timestamp 0
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_357
timestamp 0
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_363
timestamp 0
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_365
timestamp 0
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_377
timestamp 0
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_389
timestamp 0
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_401
timestamp 0
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_413
timestamp 0
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_419
timestamp 0
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_421
timestamp 0
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_433
timestamp 0
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_445
timestamp 0
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_457
timestamp 0
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_469
timestamp 0
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_475
timestamp 0
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_477
timestamp 0
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_489
timestamp 0
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_501
timestamp 0
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_513
timestamp 0
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_525
timestamp 0
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_531
timestamp 0
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_533
timestamp 0
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_545
timestamp 0
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_557
timestamp 0
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_569
timestamp 0
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_581
timestamp 0
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_587
timestamp 0
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_589
timestamp 0
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_601
timestamp 0
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_613
timestamp 0
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 0
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 0
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 0
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 0
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 0
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 0
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 0
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 0
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_81
timestamp 0
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_93
timestamp 0
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_105
timestamp 0
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 0
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 0
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_125
timestamp 0
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_137
timestamp 0
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_149
timestamp 0
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_161
timestamp 0
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 0
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 0
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_181
timestamp 0
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_193
timestamp 0
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_205
timestamp 0
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_217
timestamp 0
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 0
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 0
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_237
timestamp 0
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_249
timestamp 0
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_261
timestamp 0
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_273
timestamp 0
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 0
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 0
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_293
timestamp 0
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_305
timestamp 0
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_317
timestamp 0
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_329
timestamp 0
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_335
timestamp 0
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_337
timestamp 0
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_349
timestamp 0
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_361
timestamp 0
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_373
timestamp 0
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_385
timestamp 0
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_391
timestamp 0
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_393
timestamp 0
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_405
timestamp 0
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_417
timestamp 0
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_429
timestamp 0
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_441
timestamp 0
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_447
timestamp 0
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_449
timestamp 0
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_461
timestamp 0
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_473
timestamp 0
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_485
timestamp 0
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_497
timestamp 0
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_503
timestamp 0
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_505
timestamp 0
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_517
timestamp 0
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_529
timestamp 0
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_541
timestamp 0
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_553
timestamp 0
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_559
timestamp 0
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_561
timestamp 0
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_573
timestamp 0
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_585
timestamp 0
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_597
timestamp 0
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_609
timestamp 0
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_615
timestamp 0
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_617
timestamp 0
transform 1 0 57868 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 0
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 0
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 0
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 0
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 0
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 0
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 0
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 0
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 0
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 0
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_97
timestamp 0
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_109
timestamp 0
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_121
timestamp 0
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_133
timestamp 0
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 0
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 0
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_153
timestamp 0
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_165
timestamp 0
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_177
timestamp 0
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_189
timestamp 0
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 0
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 0
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_209
timestamp 0
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_221
timestamp 0
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_233
timestamp 0
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_245
timestamp 0
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 0
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 0
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_265
timestamp 0
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_277
timestamp 0
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_289
timestamp 0
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_301
timestamp 0
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_307
timestamp 0
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 0
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_321
timestamp 0
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_333
timestamp 0
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_345
timestamp 0
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_357
timestamp 0
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_363
timestamp 0
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_365
timestamp 0
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_377
timestamp 0
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_389
timestamp 0
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_401
timestamp 0
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_413
timestamp 0
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_419
timestamp 0
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_421
timestamp 0
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_433
timestamp 0
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_445
timestamp 0
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_457
timestamp 0
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_469
timestamp 0
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_475
timestamp 0
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_477
timestamp 0
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_489
timestamp 0
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_501
timestamp 0
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_513
timestamp 0
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_525
timestamp 0
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_531
timestamp 0
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_533
timestamp 0
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_545
timestamp 0
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_557
timestamp 0
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_569
timestamp 0
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_581
timestamp 0
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_587
timestamp 0
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_589
timestamp 0
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_601
timestamp 0
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_613
timestamp 0
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 0
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 0
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 0
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 0
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 0
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 0
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 0
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 0
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_81
timestamp 0
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_93
timestamp 0
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_105
timestamp 0
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 0
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 0
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 0
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_137
timestamp 0
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_149
timestamp 0
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 0
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 0
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 0
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 0
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_193
timestamp 0
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_205
timestamp 0
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_217
timestamp 0
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 0
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 0
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_237
timestamp 0
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_249
timestamp 0
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_261
timestamp 0
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_273
timestamp 0
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 0
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 0
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_293
timestamp 0
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_305
timestamp 0
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_317
timestamp 0
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_329
timestamp 0
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_335
timestamp 0
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_337
timestamp 0
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_349
timestamp 0
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_361
timestamp 0
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_373
timestamp 0
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_385
timestamp 0
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_391
timestamp 0
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_393
timestamp 0
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_405
timestamp 0
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_417
timestamp 0
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_429
timestamp 0
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_441
timestamp 0
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_447
timestamp 0
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_449
timestamp 0
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_461
timestamp 0
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_473
timestamp 0
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_485
timestamp 0
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_497
timestamp 0
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_503
timestamp 0
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_505
timestamp 0
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_517
timestamp 0
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_529
timestamp 0
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_541
timestamp 0
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_553
timestamp 0
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_559
timestamp 0
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_561
timestamp 0
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_573
timestamp 0
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_585
timestamp 0
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_597
timestamp 0
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_609
timestamp 0
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_615
timestamp 0
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_617
timestamp 0
transform 1 0 57868 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 0
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 0
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 0
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 0
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 0
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 0
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 0
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 0
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 0
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 0
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 0
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 0
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_121
timestamp 0
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_133
timestamp 0
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 0
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 0
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_153
timestamp 0
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_165
timestamp 0
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_177
timestamp 0
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_189
timestamp 0
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 0
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 0
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_209
timestamp 0
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_221
timestamp 0
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_233
timestamp 0
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_245
timestamp 0
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 0
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 0
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_265
timestamp 0
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_277
timestamp 0
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_289
timestamp 0
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_301
timestamp 0
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_307
timestamp 0
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 0
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_321
timestamp 0
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_333
timestamp 0
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_345
timestamp 0
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_357
timestamp 0
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_363
timestamp 0
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_365
timestamp 0
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_377
timestamp 0
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_389
timestamp 0
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_401
timestamp 0
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_413
timestamp 0
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_419
timestamp 0
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_421
timestamp 0
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_433
timestamp 0
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_445
timestamp 0
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_457
timestamp 0
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_469
timestamp 0
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_475
timestamp 0
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_477
timestamp 0
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_489
timestamp 0
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_501
timestamp 0
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_513
timestamp 0
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_525
timestamp 0
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_531
timestamp 0
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_533
timestamp 0
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_545
timestamp 0
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_557
timestamp 0
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_569
timestamp 0
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_581
timestamp 0
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_587
timestamp 0
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_589
timestamp 0
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_601
timestamp 0
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_613
timestamp 0
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 0
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 0
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 0
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 0
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 0
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 0
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 0
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 0
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 0
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 0
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_105
timestamp 0
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 0
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 0
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_125
timestamp 0
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_137
timestamp 0
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_149
timestamp 0
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_161
timestamp 0
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 0
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 0
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_181
timestamp 0
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_193
timestamp 0
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_205
timestamp 0
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_217
timestamp 0
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 0
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 0
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 0
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 0
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_261
timestamp 0
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_273
timestamp 0
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 0
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 0
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_293
timestamp 0
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_305
timestamp 0
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_317
timestamp 0
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_329
timestamp 0
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_335
timestamp 0
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 0
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_349
timestamp 0
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_361
timestamp 0
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_373
timestamp 0
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_385
timestamp 0
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_391
timestamp 0
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_393
timestamp 0
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_405
timestamp 0
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_417
timestamp 0
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_429
timestamp 0
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_441
timestamp 0
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_447
timestamp 0
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_449
timestamp 0
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_461
timestamp 0
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_473
timestamp 0
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_485
timestamp 0
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_497
timestamp 0
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_503
timestamp 0
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_505
timestamp 0
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_517
timestamp 0
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_529
timestamp 0
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_541
timestamp 0
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_553
timestamp 0
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_559
timestamp 0
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_561
timestamp 0
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_573
timestamp 0
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_585
timestamp 0
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_597
timestamp 0
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_609
timestamp 0
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_615
timestamp 0
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_617
timestamp 0
transform 1 0 57868 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 0
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 0
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 0
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 0
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 0
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 0
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 0
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 0
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 0
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 0
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 0
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_109
timestamp 0
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_121
timestamp 0
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_133
timestamp 0
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 0
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 0
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_153
timestamp 0
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_165
timestamp 0
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_177
timestamp 0
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_189
timestamp 0
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 0
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_197
timestamp 0
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_209
timestamp 0
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_221
timestamp 0
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_233
timestamp 0
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_245
timestamp 0
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 0
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 0
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 0
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_277
timestamp 0
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_289
timestamp 0
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_301
timestamp 0
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_307
timestamp 0
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_309
timestamp 0
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_321
timestamp 0
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_333
timestamp 0
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_345
timestamp 0
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_357
timestamp 0
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_363
timestamp 0
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_365
timestamp 0
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_377
timestamp 0
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_389
timestamp 0
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_401
timestamp 0
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_413
timestamp 0
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_419
timestamp 0
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_421
timestamp 0
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_433
timestamp 0
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_445
timestamp 0
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_457
timestamp 0
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_469
timestamp 0
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_475
timestamp 0
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_477
timestamp 0
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_489
timestamp 0
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_501
timestamp 0
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_513
timestamp 0
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_525
timestamp 0
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_531
timestamp 0
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_533
timestamp 0
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_545
timestamp 0
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_557
timestamp 0
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_569
timestamp 0
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_581
timestamp 0
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_587
timestamp 0
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_589
timestamp 0
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_601
timestamp 0
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_613
timestamp 0
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 0
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 0
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 0
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 0
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 0
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 0
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 0
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 0
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 0
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_93
timestamp 0
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_105
timestamp 0
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 0
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 0
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 0
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 0
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 0
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 0
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 0
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 0
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_181
timestamp 0
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_193
timestamp 0
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_205
timestamp 0
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_217
timestamp 0
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 0
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 0
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 0
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_249
timestamp 0
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_261
timestamp 0
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_273
timestamp 0
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 0
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 0
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 0
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_305
timestamp 0
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_317
timestamp 0
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_329
timestamp 0
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_335
timestamp 0
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_337
timestamp 0
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_349
timestamp 0
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_361
timestamp 0
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_373
timestamp 0
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_385
timestamp 0
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_391
timestamp 0
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_393
timestamp 0
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_405
timestamp 0
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_417
timestamp 0
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_429
timestamp 0
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_441
timestamp 0
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_447
timestamp 0
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_449
timestamp 0
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_461
timestamp 0
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_473
timestamp 0
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_485
timestamp 0
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_497
timestamp 0
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_503
timestamp 0
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_505
timestamp 0
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_517
timestamp 0
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_529
timestamp 0
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_541
timestamp 0
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_553
timestamp 0
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_559
timestamp 0
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_561
timestamp 0
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_573
timestamp 0
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_585
timestamp 0
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_597
timestamp 0
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_609
timestamp 0
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_615
timestamp 0
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_617
timestamp 0
transform 1 0 57868 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 0
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 0
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 0
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 0
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 0
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 0
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 0
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 0
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 0
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 0
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 0
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_109
timestamp 0
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_121
timestamp 0
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_133
timestamp 0
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 0
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 0
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 0
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_165
timestamp 0
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_177
timestamp 0
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_189
timestamp 0
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 0
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 0
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_209
timestamp 0
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_221
timestamp 0
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_233
timestamp 0
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_245
timestamp 0
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 0
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 0
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 0
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 0
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_289
timestamp 0
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_301
timestamp 0
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 0
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_309
timestamp 0
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_321
timestamp 0
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_333
timestamp 0
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_345
timestamp 0
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_357
timestamp 0
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_363
timestamp 0
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_365
timestamp 0
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_377
timestamp 0
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_389
timestamp 0
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_401
timestamp 0
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_413
timestamp 0
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_419
timestamp 0
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_421
timestamp 0
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_433
timestamp 0
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_445
timestamp 0
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_457
timestamp 0
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_469
timestamp 0
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_475
timestamp 0
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_477
timestamp 0
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_489
timestamp 0
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_501
timestamp 0
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_513
timestamp 0
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_525
timestamp 0
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_531
timestamp 0
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_533
timestamp 0
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_545
timestamp 0
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_557
timestamp 0
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_569
timestamp 0
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_581
timestamp 0
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_587
timestamp 0
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_589
timestamp 0
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_601
timestamp 0
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_613
timestamp 0
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 0
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 0
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 0
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 0
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 0
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 0
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 0
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 0
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 0
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 0
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 0
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 0
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 0
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 0
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_137
timestamp 0
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_149
timestamp 0
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_161
timestamp 0
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 0
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 0
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_181
timestamp 0
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_193
timestamp 0
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_205
timestamp 0
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_217
timestamp 0
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 0
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 0
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 0
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 0
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 0
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_273
timestamp 0
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 0
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 0
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_293
timestamp 0
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_305
timestamp 0
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_317
timestamp 0
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_329
timestamp 0
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 0
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_337
timestamp 0
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_349
timestamp 0
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_361
timestamp 0
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_373
timestamp 0
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_385
timestamp 0
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_391
timestamp 0
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_393
timestamp 0
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_405
timestamp 0
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_417
timestamp 0
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_429
timestamp 0
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_441
timestamp 0
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_447
timestamp 0
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_449
timestamp 0
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_461
timestamp 0
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_473
timestamp 0
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_485
timestamp 0
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_497
timestamp 0
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_503
timestamp 0
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_505
timestamp 0
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_517
timestamp 0
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_529
timestamp 0
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_541
timestamp 0
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_553
timestamp 0
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_559
timestamp 0
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_561
timestamp 0
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_573
timestamp 0
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_585
timestamp 0
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_597
timestamp 0
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_609
timestamp 0
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_615
timestamp 0
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_617
timestamp 0
transform 1 0 57868 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 0
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 0
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 0
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 0
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 0
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 0
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_65
timestamp 0
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_77
timestamp 0
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 0
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 0
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 0
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 0
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_121
timestamp 0
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 0
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 0
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 0
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_153
timestamp 0
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_165
timestamp 0
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_177
timestamp 0
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_189
timestamp 0
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 0
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 0
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 0
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_221
timestamp 0
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_233
timestamp 0
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_245
timestamp 0
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 0
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 0
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 0
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_277
timestamp 0
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_289
timestamp 0
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_301
timestamp 0
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_307
timestamp 0
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 0
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_321
timestamp 0
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_333
timestamp 0
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_345
timestamp 0
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_357
timestamp 0
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_363
timestamp 0
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_365
timestamp 0
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_377
timestamp 0
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_389
timestamp 0
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_401
timestamp 0
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_413
timestamp 0
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_419
timestamp 0
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_421
timestamp 0
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_433
timestamp 0
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_445
timestamp 0
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_457
timestamp 0
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_469
timestamp 0
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_475
timestamp 0
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_477
timestamp 0
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_489
timestamp 0
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_501
timestamp 0
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_513
timestamp 0
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_525
timestamp 0
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_531
timestamp 0
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_533
timestamp 0
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_545
timestamp 0
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_557
timestamp 0
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_569
timestamp 0
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_581
timestamp 0
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_587
timestamp 0
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_589
timestamp 0
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_601
timestamp 0
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_613
timestamp 0
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 0
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 0
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 0
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 0
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 0
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 0
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 0
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 0
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_81
timestamp 0
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_93
timestamp 0
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_105
timestamp 0
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 0
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 0
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_125
timestamp 0
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_137
timestamp 0
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_149
timestamp 0
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_161
timestamp 0
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 0
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 0
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_181
timestamp 0
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_193
timestamp 0
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_205
timestamp 0
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_217
timestamp 0
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 0
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_225
timestamp 0
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_237
timestamp 0
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_249
timestamp 0
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_261
timestamp 0
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_273
timestamp 0
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 0
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 0
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 0
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 0
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_317
timestamp 0
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_329
timestamp 0
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_335
timestamp 0
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_337
timestamp 0
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_349
timestamp 0
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_361
timestamp 0
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_373
timestamp 0
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_385
timestamp 0
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_391
timestamp 0
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_393
timestamp 0
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_405
timestamp 0
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_417
timestamp 0
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_429
timestamp 0
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_441
timestamp 0
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_447
timestamp 0
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_449
timestamp 0
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_461
timestamp 0
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_473
timestamp 0
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_485
timestamp 0
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_497
timestamp 0
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_503
timestamp 0
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_505
timestamp 0
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_517
timestamp 0
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_529
timestamp 0
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_541
timestamp 0
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_553
timestamp 0
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_559
timestamp 0
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_561
timestamp 0
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_573
timestamp 0
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_585
timestamp 0
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_597
timestamp 0
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_609
timestamp 0
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_615
timestamp 0
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_617
timestamp 0
transform 1 0 57868 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 0
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 0
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 0
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 0
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 0
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 0
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 0
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_77
timestamp 0
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 0
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 0
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_97
timestamp 0
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_109
timestamp 0
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_121
timestamp 0
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_133
timestamp 0
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 0
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 0
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 0
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_165
timestamp 0
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_177
timestamp 0
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_189
timestamp 0
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 0
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_197
timestamp 0
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_209
timestamp 0
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_221
timestamp 0
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_233
timestamp 0
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_245
timestamp 0
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 0
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 0
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 0
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_277
timestamp 0
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_289
timestamp 0
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_301
timestamp 0
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 0
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 0
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_321
timestamp 0
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_333
timestamp 0
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_345
timestamp 0
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_357
timestamp 0
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_363
timestamp 0
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_365
timestamp 0
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_377
timestamp 0
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_389
timestamp 0
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_401
timestamp 0
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_413
timestamp 0
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_419
timestamp 0
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_421
timestamp 0
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_433
timestamp 0
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_445
timestamp 0
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_457
timestamp 0
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_469
timestamp 0
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_475
timestamp 0
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_477
timestamp 0
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_489
timestamp 0
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_501
timestamp 0
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_513
timestamp 0
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_525
timestamp 0
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_531
timestamp 0
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_533
timestamp 0
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_545
timestamp 0
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_557
timestamp 0
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_569
timestamp 0
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_581
timestamp 0
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_587
timestamp 0
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_589
timestamp 0
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_601
timestamp 0
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_613
timestamp 0
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 0
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 0
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 0
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_39
timestamp 0
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 0
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 0
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 0
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 0
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_81
timestamp 0
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_93
timestamp 0
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_105
timestamp 0
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_111
timestamp 0
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 0
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_125
timestamp 0
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_137
timestamp 0
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_149
timestamp 0
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_161
timestamp 0
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 0
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 0
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_181
timestamp 0
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_193
timestamp 0
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_205
timestamp 0
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_217
timestamp 0
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_223
timestamp 0
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_225
timestamp 0
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_237
timestamp 0
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_249
timestamp 0
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_261
timestamp 0
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_273
timestamp 0
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 0
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 0
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 0
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_305
timestamp 0
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_317
timestamp 0
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_329
timestamp 0
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_335
timestamp 0
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_337
timestamp 0
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_349
timestamp 0
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_361
timestamp 0
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_373
timestamp 0
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_385
timestamp 0
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_391
timestamp 0
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_393
timestamp 0
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_405
timestamp 0
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_417
timestamp 0
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_429
timestamp 0
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_441
timestamp 0
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_447
timestamp 0
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_449
timestamp 0
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_461
timestamp 0
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_473
timestamp 0
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_485
timestamp 0
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_497
timestamp 0
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_503
timestamp 0
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_505
timestamp 0
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_517
timestamp 0
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_529
timestamp 0
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_541
timestamp 0
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_553
timestamp 0
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_559
timestamp 0
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_561
timestamp 0
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_573
timestamp 0
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_585
timestamp 0
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_597
timestamp 0
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_609
timestamp 0
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_615
timestamp 0
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_617
timestamp 0
transform 1 0 57868 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 0
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 0
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 0
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 0
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 0
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 0
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_65
timestamp 0
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 0
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 0
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 0
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_97
timestamp 0
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_109
timestamp 0
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_121
timestamp 0
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_133
timestamp 0
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 0
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_141
timestamp 0
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_153
timestamp 0
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_165
timestamp 0
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_177
timestamp 0
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_189
timestamp 0
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 0
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 0
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_209
timestamp 0
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_221
timestamp 0
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_233
timestamp 0
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_245
timestamp 0
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_251
timestamp 0
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 0
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_265
timestamp 0
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 0
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_289
timestamp 0
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_301
timestamp 0
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 0
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 0
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_321
timestamp 0
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_333
timestamp 0
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_345
timestamp 0
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_357
timestamp 0
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_363
timestamp 0
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_365
timestamp 0
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_377
timestamp 0
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_389
timestamp 0
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_401
timestamp 0
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_413
timestamp 0
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_419
timestamp 0
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_421
timestamp 0
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_433
timestamp 0
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_445
timestamp 0
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_457
timestamp 0
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_469
timestamp 0
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_475
timestamp 0
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_477
timestamp 0
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_489
timestamp 0
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_501
timestamp 0
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_513
timestamp 0
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_525
timestamp 0
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_531
timestamp 0
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_533
timestamp 0
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_545
timestamp 0
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_557
timestamp 0
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_569
timestamp 0
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_581
timestamp 0
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_587
timestamp 0
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_589
timestamp 0
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_601
timestamp 0
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_613
timestamp 0
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 0
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 0
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 0
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 0
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 0
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 0
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 0
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 0
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 0
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_93
timestamp 0
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_105
timestamp 0
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 0
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 0
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_125
timestamp 0
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_137
timestamp 0
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 0
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_161
timestamp 0
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 0
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 0
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_181
timestamp 0
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_193
timestamp 0
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_205
timestamp 0
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_217
timestamp 0
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 0
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 0
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_237
timestamp 0
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_249
timestamp 0
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_261
timestamp 0
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_273
timestamp 0
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 0
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 0
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 0
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_305
timestamp 0
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_317
timestamp 0
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_329
timestamp 0
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 0
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_337
timestamp 0
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_349
timestamp 0
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_361
timestamp 0
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_373
timestamp 0
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_385
timestamp 0
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_391
timestamp 0
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_393
timestamp 0
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_405
timestamp 0
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_417
timestamp 0
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_429
timestamp 0
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_441
timestamp 0
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_447
timestamp 0
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_449
timestamp 0
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_461
timestamp 0
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_473
timestamp 0
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_485
timestamp 0
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_497
timestamp 0
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_503
timestamp 0
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_505
timestamp 0
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_517
timestamp 0
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_529
timestamp 0
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_541
timestamp 0
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_553
timestamp 0
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_559
timestamp 0
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_561
timestamp 0
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_573
timestamp 0
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_585
timestamp 0
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_597
timestamp 0
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_609
timestamp 0
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_615
timestamp 0
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_617
timestamp 0
transform 1 0 57868 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 0
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 0
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 0
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 0
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 0
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 0
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 0
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 0
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 0
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 0
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_97
timestamp 0
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_109
timestamp 0
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_121
timestamp 0
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_133
timestamp 0
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 0
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 0
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_153
timestamp 0
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_165
timestamp 0
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_177
timestamp 0
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_189
timestamp 0
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_195
timestamp 0
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 0
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_209
timestamp 0
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_221
timestamp 0
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_233
timestamp 0
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_245
timestamp 0
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 0
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_253
timestamp 0
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_265
timestamp 0
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_277
timestamp 0
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_289
timestamp 0
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_301
timestamp 0
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 0
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 0
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_321
timestamp 0
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_333
timestamp 0
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_345
timestamp 0
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_357
timestamp 0
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_363
timestamp 0
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_365
timestamp 0
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_377
timestamp 0
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_389
timestamp 0
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_401
timestamp 0
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_413
timestamp 0
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_419
timestamp 0
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_421
timestamp 0
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_433
timestamp 0
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_445
timestamp 0
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_457
timestamp 0
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_469
timestamp 0
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_475
timestamp 0
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_477
timestamp 0
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_489
timestamp 0
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_501
timestamp 0
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_513
timestamp 0
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_525
timestamp 0
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_531
timestamp 0
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_533
timestamp 0
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_545
timestamp 0
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_557
timestamp 0
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_569
timestamp 0
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_581
timestamp 0
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_587
timestamp 0
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_589
timestamp 0
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_601
timestamp 0
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_613
timestamp 0
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 0
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 0
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 0
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 0
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 0
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 0
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 0
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 0
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_81
timestamp 0
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_93
timestamp 0
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_105
timestamp 0
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 0
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 0
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 0
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_137
timestamp 0
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_149
timestamp 0
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_161
timestamp 0
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 0
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 0
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_181
timestamp 0
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_193
timestamp 0
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_205
timestamp 0
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_217
timestamp 0
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 0
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_225
timestamp 0
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_237
timestamp 0
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_249
timestamp 0
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_261
timestamp 0
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_273
timestamp 0
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 0
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_281
timestamp 0
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_293
timestamp 0
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_305
timestamp 0
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_317
timestamp 0
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_329
timestamp 0
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 0
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_337
timestamp 0
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_349
timestamp 0
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_361
timestamp 0
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_373
timestamp 0
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_385
timestamp 0
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_391
timestamp 0
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_393
timestamp 0
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_405
timestamp 0
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_417
timestamp 0
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_429
timestamp 0
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_441
timestamp 0
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_447
timestamp 0
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_449
timestamp 0
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_461
timestamp 0
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_473
timestamp 0
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_485
timestamp 0
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_497
timestamp 0
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_503
timestamp 0
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_505
timestamp 0
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_517
timestamp 0
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_529
timestamp 0
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_541
timestamp 0
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_553
timestamp 0
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_559
timestamp 0
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_561
timestamp 0
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_573
timestamp 0
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_585
timestamp 0
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_597
timestamp 0
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_609
timestamp 0
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_615
timestamp 0
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_617
timestamp 0
transform 1 0 57868 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 0
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 0
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 0
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 0
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 0
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 0
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 0
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 0
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 0
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 0
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_97
timestamp 0
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_109
timestamp 0
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_121
timestamp 0
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_133
timestamp 0
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 0
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 0
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 0
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_165
timestamp 0
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_177
timestamp 0
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_189
timestamp 0
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 0
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_197
timestamp 0
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_209
timestamp 0
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_221
timestamp 0
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_233
timestamp 0
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_245
timestamp 0
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_251
timestamp 0
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_253
timestamp 0
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_265
timestamp 0
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_277
timestamp 0
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_289
timestamp 0
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_301
timestamp 0
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_307
timestamp 0
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_309
timestamp 0
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_321
timestamp 0
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_333
timestamp 0
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_345
timestamp 0
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_357
timestamp 0
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_363
timestamp 0
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_365
timestamp 0
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_377
timestamp 0
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_389
timestamp 0
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_401
timestamp 0
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_413
timestamp 0
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_419
timestamp 0
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_421
timestamp 0
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_433
timestamp 0
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_445
timestamp 0
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_457
timestamp 0
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_469
timestamp 0
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_475
timestamp 0
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_477
timestamp 0
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_489
timestamp 0
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_501
timestamp 0
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_513
timestamp 0
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_525
timestamp 0
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_531
timestamp 0
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_533
timestamp 0
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_545
timestamp 0
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_557
timestamp 0
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_569
timestamp 0
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_581
timestamp 0
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_587
timestamp 0
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_589
timestamp 0
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_601
timestamp 0
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_613
timestamp 0
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 0
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 0
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 0
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 0
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_51
timestamp 0
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 0
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 0
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 0
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 0
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_93
timestamp 0
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_105
timestamp 0
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 0
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 0
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_125
timestamp 0
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_137
timestamp 0
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_149
timestamp 0
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_161
timestamp 0
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 0
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 0
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_181
timestamp 0
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_193
timestamp 0
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_205
timestamp 0
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_217
timestamp 0
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 0
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 0
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_237
timestamp 0
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_249
timestamp 0
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_261
timestamp 0
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_273
timestamp 0
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 0
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_281
timestamp 0
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_293
timestamp 0
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_305
timestamp 0
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_317
timestamp 0
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_329
timestamp 0
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 0
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_337
timestamp 0
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_349
timestamp 0
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_361
timestamp 0
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_373
timestamp 0
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_385
timestamp 0
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_391
timestamp 0
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_393
timestamp 0
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_405
timestamp 0
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_417
timestamp 0
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_429
timestamp 0
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_441
timestamp 0
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_447
timestamp 0
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_449
timestamp 0
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_461
timestamp 0
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_473
timestamp 0
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_485
timestamp 0
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_497
timestamp 0
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_503
timestamp 0
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_505
timestamp 0
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_517
timestamp 0
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_529
timestamp 0
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_541
timestamp 0
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_553
timestamp 0
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_559
timestamp 0
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_561
timestamp 0
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_573
timestamp 0
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_585
timestamp 0
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_597
timestamp 0
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_609
timestamp 0
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_615
timestamp 0
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_617
timestamp 0
transform 1 0 57868 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 0
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 0
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 0
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 0
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 0
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 0
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_65
timestamp 0
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 0
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 0
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 0
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 0
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 0
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 0
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 0
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 0
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 0
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 0
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_165
timestamp 0
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_177
timestamp 0
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_189
timestamp 0
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 0
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 0
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_209
timestamp 0
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_221
timestamp 0
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_233
timestamp 0
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 0
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 0
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 0
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_265
timestamp 0
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_277
timestamp 0
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_289
timestamp 0
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_301
timestamp 0
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 0
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_309
timestamp 0
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_321
timestamp 0
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_333
timestamp 0
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_345
timestamp 0
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_357
timestamp 0
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_363
timestamp 0
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_365
timestamp 0
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_377
timestamp 0
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_389
timestamp 0
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_401
timestamp 0
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_413
timestamp 0
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_419
timestamp 0
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_421
timestamp 0
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_433
timestamp 0
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_445
timestamp 0
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_457
timestamp 0
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_469
timestamp 0
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_475
timestamp 0
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_477
timestamp 0
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_489
timestamp 0
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_501
timestamp 0
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_513
timestamp 0
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_525
timestamp 0
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_531
timestamp 0
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_533
timestamp 0
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_545
timestamp 0
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_557
timestamp 0
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_569
timestamp 0
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_581
timestamp 0
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_587
timestamp 0
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_589
timestamp 0
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_601
timestamp 0
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_613
timestamp 0
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 0
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 0
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 0
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 0
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 0
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 0
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 0
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_69
timestamp 0
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_81
timestamp 0
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_93
timestamp 0
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_105
timestamp 0
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 0
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 0
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 0
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_137
timestamp 0
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_149
timestamp 0
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_161
timestamp 0
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 0
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 0
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_181
timestamp 0
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_193
timestamp 0
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_205
timestamp 0
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_217
timestamp 0
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_223
timestamp 0
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_225
timestamp 0
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_237
timestamp 0
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_249
timestamp 0
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_261
timestamp 0
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_273
timestamp 0
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_279
timestamp 0
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_281
timestamp 0
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_293
timestamp 0
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_305
timestamp 0
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_317
timestamp 0
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_329
timestamp 0
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_335
timestamp 0
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_337
timestamp 0
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_349
timestamp 0
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_361
timestamp 0
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_373
timestamp 0
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_385
timestamp 0
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_391
timestamp 0
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_393
timestamp 0
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_405
timestamp 0
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_417
timestamp 0
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_429
timestamp 0
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_441
timestamp 0
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_447
timestamp 0
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_449
timestamp 0
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_461
timestamp 0
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_473
timestamp 0
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_485
timestamp 0
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_497
timestamp 0
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_503
timestamp 0
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_505
timestamp 0
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_517
timestamp 0
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_529
timestamp 0
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_541
timestamp 0
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_553
timestamp 0
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_559
timestamp 0
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_561
timestamp 0
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_573
timestamp 0
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_585
timestamp 0
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_597
timestamp 0
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_609
timestamp 0
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_615
timestamp 0
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_617
timestamp 0
transform 1 0 57868 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 0
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 0
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 0
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 0
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 0
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 0
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 0
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 0
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 0
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 0
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 0
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_109
timestamp 0
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_121
timestamp 0
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_133
timestamp 0
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 0
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_141
timestamp 0
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_153
timestamp 0
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_165
timestamp 0
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_177
timestamp 0
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_189
timestamp 0
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 0
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 0
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_209
timestamp 0
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_221
timestamp 0
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_233
timestamp 0
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_245
timestamp 0
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_251
timestamp 0
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_253
timestamp 0
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_265
timestamp 0
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_277
timestamp 0
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_289
timestamp 0
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_301
timestamp 0
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_307
timestamp 0
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_309
timestamp 0
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_321
timestamp 0
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_333
timestamp 0
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_345
timestamp 0
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_357
timestamp 0
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_363
timestamp 0
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_365
timestamp 0
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_377
timestamp 0
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_389
timestamp 0
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_401
timestamp 0
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_413
timestamp 0
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_419
timestamp 0
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_421
timestamp 0
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_433
timestamp 0
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_445
timestamp 0
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_457
timestamp 0
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_469
timestamp 0
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_475
timestamp 0
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_477
timestamp 0
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_489
timestamp 0
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_501
timestamp 0
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_513
timestamp 0
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_525
timestamp 0
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_531
timestamp 0
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_533
timestamp 0
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_545
timestamp 0
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_557
timestamp 0
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_569
timestamp 0
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_581
timestamp 0
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_587
timestamp 0
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_589
timestamp 0
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_601
timestamp 0
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_613
timestamp 0
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 0
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 0
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 0
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 0
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 0
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 0
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 0
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 0
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 0
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_93
timestamp 0
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_105
timestamp 0
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 0
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_113
timestamp 0
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_125
timestamp 0
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_137
timestamp 0
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_149
timestamp 0
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_161
timestamp 0
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 0
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 0
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_181
timestamp 0
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_193
timestamp 0
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_205
timestamp 0
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_217
timestamp 0
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_223
timestamp 0
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_225
timestamp 0
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_237
timestamp 0
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_249
timestamp 0
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_261
timestamp 0
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_273
timestamp 0
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 0
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 0
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_293
timestamp 0
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_305
timestamp 0
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_317
timestamp 0
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_329
timestamp 0
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 0
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 0
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 0
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_361
timestamp 0
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_373
timestamp 0
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_385
timestamp 0
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_391
timestamp 0
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_393
timestamp 0
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_405
timestamp 0
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_417
timestamp 0
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_429
timestamp 0
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_441
timestamp 0
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_447
timestamp 0
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_449
timestamp 0
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_461
timestamp 0
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_473
timestamp 0
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_485
timestamp 0
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_497
timestamp 0
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_503
timestamp 0
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_505
timestamp 0
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_517
timestamp 0
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_529
timestamp 0
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_541
timestamp 0
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_553
timestamp 0
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_559
timestamp 0
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_561
timestamp 0
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_573
timestamp 0
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_585
timestamp 0
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_597
timestamp 0
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_609
timestamp 0
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_615
timestamp 0
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_617
timestamp 0
transform 1 0 57868 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 0
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 0
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 0
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 0
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 0
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 0
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 0
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 0
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 0
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_85
timestamp 0
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_97
timestamp 0
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_109
timestamp 0
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_121
timestamp 0
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_133
timestamp 0
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 0
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 0
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 0
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_165
timestamp 0
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_177
timestamp 0
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_189
timestamp 0
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 0
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 0
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 0
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_221
timestamp 0
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_233
timestamp 0
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_245
timestamp 0
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_251
timestamp 0
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_253
timestamp 0
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_265
timestamp 0
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_277
timestamp 0
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_289
timestamp 0
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_301
timestamp 0
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 0
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 0
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 0
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_333
timestamp 0
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_345
timestamp 0
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_357
timestamp 0
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 0
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_365
timestamp 0
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_377
timestamp 0
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_389
timestamp 0
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_401
timestamp 0
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_413
timestamp 0
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_419
timestamp 0
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_421
timestamp 0
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_433
timestamp 0
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_445
timestamp 0
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_457
timestamp 0
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_469
timestamp 0
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_475
timestamp 0
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_477
timestamp 0
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_489
timestamp 0
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_501
timestamp 0
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_513
timestamp 0
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_525
timestamp 0
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_531
timestamp 0
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_533
timestamp 0
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_545
timestamp 0
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_557
timestamp 0
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_569
timestamp 0
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_581
timestamp 0
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_587
timestamp 0
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_589
timestamp 0
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_601
timestamp 0
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_613
timestamp 0
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 0
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 0
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 0
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 0
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 0
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 0
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 0
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 0
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_81
timestamp 0
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_93
timestamp 0
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_105
timestamp 0
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 0
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 0
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 0
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_137
timestamp 0
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_149
timestamp 0
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_161
timestamp 0
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 0
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 0
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 0
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_193
timestamp 0
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_205
timestamp 0
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_217
timestamp 0
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 0
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_225
timestamp 0
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_237
timestamp 0
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_249
timestamp 0
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_261
timestamp 0
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_273
timestamp 0
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 0
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 0
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 0
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_305
timestamp 0
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_317
timestamp 0
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_329
timestamp 0
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_335
timestamp 0
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 0
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 0
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_361
timestamp 0
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_373
timestamp 0
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_385
timestamp 0
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_391
timestamp 0
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_393
timestamp 0
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_405
timestamp 0
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_417
timestamp 0
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_429
timestamp 0
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_441
timestamp 0
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_447
timestamp 0
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_449
timestamp 0
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_461
timestamp 0
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_473
timestamp 0
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_485
timestamp 0
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_497
timestamp 0
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_503
timestamp 0
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_505
timestamp 0
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_517
timestamp 0
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_529
timestamp 0
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_541
timestamp 0
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_553
timestamp 0
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_559
timestamp 0
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_561
timestamp 0
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_573
timestamp 0
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_585
timestamp 0
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_597
timestamp 0
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_609
timestamp 0
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_615
timestamp 0
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_617
timestamp 0
transform 1 0 57868 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 0
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 0
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 0
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 0
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 0
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 0
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_65
timestamp 0
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_77
timestamp 0
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 0
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_85
timestamp 0
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_97
timestamp 0
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_109
timestamp 0
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_121
timestamp 0
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_133
timestamp 0
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_139
timestamp 0
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 0
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_153
timestamp 0
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_165
timestamp 0
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_177
timestamp 0
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_189
timestamp 0
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_195
timestamp 0
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_197
timestamp 0
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_209
timestamp 0
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_221
timestamp 0
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_233
timestamp 0
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_245
timestamp 0
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_251
timestamp 0
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 0
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_265
timestamp 0
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_277
timestamp 0
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_289
timestamp 0
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_301
timestamp 0
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_307
timestamp 0
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 0
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 0
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_333
timestamp 0
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_345
timestamp 0
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_357
timestamp 0
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_363
timestamp 0
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_365
timestamp 0
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_377
timestamp 0
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_389
timestamp 0
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_401
timestamp 0
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_413
timestamp 0
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_419
timestamp 0
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_421
timestamp 0
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_433
timestamp 0
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_445
timestamp 0
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_457
timestamp 0
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_469
timestamp 0
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_475
timestamp 0
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_477
timestamp 0
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_489
timestamp 0
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_501
timestamp 0
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_513
timestamp 0
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_525
timestamp 0
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_531
timestamp 0
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_533
timestamp 0
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_545
timestamp 0
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_557
timestamp 0
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_569
timestamp 0
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_581
timestamp 0
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_587
timestamp 0
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_589
timestamp 0
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_601
timestamp 0
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_613
timestamp 0
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 0
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 0
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 0
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 0
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 0
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 0
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 0
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 0
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_81
timestamp 0
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_93
timestamp 0
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_105
timestamp 0
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_111
timestamp 0
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_113
timestamp 0
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_125
timestamp 0
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_137
timestamp 0
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_149
timestamp 0
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_161
timestamp 0
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_167
timestamp 0
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_169
timestamp 0
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_181
timestamp 0
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_193
timestamp 0
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_205
timestamp 0
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_217
timestamp 0
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_223
timestamp 0
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_225
timestamp 0
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_237
timestamp 0
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_249
timestamp 0
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_261
timestamp 0
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_273
timestamp 0
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_279
timestamp 0
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_281
timestamp 0
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_293
timestamp 0
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_305
timestamp 0
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_317
timestamp 0
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_329
timestamp 0
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_335
timestamp 0
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_337
timestamp 0
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_349
timestamp 0
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_361
timestamp 0
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_373
timestamp 0
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_385
timestamp 0
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_391
timestamp 0
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_393
timestamp 0
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_405
timestamp 0
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_417
timestamp 0
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_429
timestamp 0
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_441
timestamp 0
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_447
timestamp 0
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_449
timestamp 0
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_461
timestamp 0
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_473
timestamp 0
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_485
timestamp 0
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_497
timestamp 0
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_503
timestamp 0
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_505
timestamp 0
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_517
timestamp 0
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_529
timestamp 0
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_541
timestamp 0
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_553
timestamp 0
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_559
timestamp 0
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_561
timestamp 0
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_573
timestamp 0
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_585
timestamp 0
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_597
timestamp 0
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_609
timestamp 0
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_615
timestamp 0
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_617
timestamp 0
transform 1 0 57868 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_3
timestamp 0
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_15
timestamp 0
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 0
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 0
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 0
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_53
timestamp 0
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_65
timestamp 0
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_77
timestamp 0
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_83
timestamp 0
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 0
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_97
timestamp 0
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_109
timestamp 0
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_121
timestamp 0
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_133
timestamp 0
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_139
timestamp 0
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 0
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_153
timestamp 0
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_165
timestamp 0
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_177
timestamp 0
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_189
timestamp 0
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_195
timestamp 0
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_197
timestamp 0
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_209
timestamp 0
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_221
timestamp 0
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_233
timestamp 0
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_245
timestamp 0
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_251
timestamp 0
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_253
timestamp 0
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_265
timestamp 0
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_277
timestamp 0
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_289
timestamp 0
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_301
timestamp 0
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_307
timestamp 0
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_309
timestamp 0
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_321
timestamp 0
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_333
timestamp 0
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_345
timestamp 0
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_357
timestamp 0
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_363
timestamp 0
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_365
timestamp 0
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_377
timestamp 0
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_389
timestamp 0
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_401
timestamp 0
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_413
timestamp 0
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_419
timestamp 0
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_421
timestamp 0
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_433
timestamp 0
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_445
timestamp 0
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_457
timestamp 0
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_469
timestamp 0
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_475
timestamp 0
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_477
timestamp 0
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_489
timestamp 0
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_501
timestamp 0
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_513
timestamp 0
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_525
timestamp 0
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_531
timestamp 0
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_533
timestamp 0
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_545
timestamp 0
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_557
timestamp 0
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_569
timestamp 0
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_581
timestamp 0
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_587
timestamp 0
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_589
timestamp 0
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_601
timestamp 0
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_613
timestamp 0
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_3
timestamp 0
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_15
timestamp 0
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_27
timestamp 0
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_39
timestamp 0
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_51
timestamp 0
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_55
timestamp 0
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_57
timestamp 0
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_69
timestamp 0
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_81
timestamp 0
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_93
timestamp 0
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_105
timestamp 0
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_111
timestamp 0
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_113
timestamp 0
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_125
timestamp 0
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_137
timestamp 0
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_149
timestamp 0
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_161
timestamp 0
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_167
timestamp 0
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_169
timestamp 0
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_181
timestamp 0
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_193
timestamp 0
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_205
timestamp 0
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_217
timestamp 0
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_223
timestamp 0
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_225
timestamp 0
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_237
timestamp 0
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_249
timestamp 0
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_261
timestamp 0
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_273
timestamp 0
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_279
timestamp 0
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_281
timestamp 0
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_293
timestamp 0
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_305
timestamp 0
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_317
timestamp 0
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_329
timestamp 0
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_335
timestamp 0
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_337
timestamp 0
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_349
timestamp 0
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_361
timestamp 0
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_373
timestamp 0
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_385
timestamp 0
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_391
timestamp 0
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_393
timestamp 0
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_405
timestamp 0
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_417
timestamp 0
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_429
timestamp 0
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_441
timestamp 0
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_447
timestamp 0
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_449
timestamp 0
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_461
timestamp 0
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_473
timestamp 0
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_485
timestamp 0
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_497
timestamp 0
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_503
timestamp 0
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_505
timestamp 0
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_517
timestamp 0
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_529
timestamp 0
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_541
timestamp 0
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_553
timestamp 0
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_559
timestamp 0
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_561
timestamp 0
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_573
timestamp 0
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_585
timestamp 0
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_597
timestamp 0
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_609
timestamp 0
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_615
timestamp 0
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_617
timestamp 0
transform 1 0 57868 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_3
timestamp 0
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_15
timestamp 0
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 0
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_29
timestamp 0
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_41
timestamp 0
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_53
timestamp 0
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_65
timestamp 0
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_77
timestamp 0
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_83
timestamp 0
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_85
timestamp 0
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_97
timestamp 0
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_109
timestamp 0
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_121
timestamp 0
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_133
timestamp 0
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_139
timestamp 0
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_141
timestamp 0
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_153
timestamp 0
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_165
timestamp 0
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_177
timestamp 0
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_189
timestamp 0
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_195
timestamp 0
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_197
timestamp 0
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_209
timestamp 0
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_221
timestamp 0
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_233
timestamp 0
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_245
timestamp 0
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_251
timestamp 0
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_253
timestamp 0
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_265
timestamp 0
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_277
timestamp 0
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_289
timestamp 0
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_301
timestamp 0
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_307
timestamp 0
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_309
timestamp 0
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_321
timestamp 0
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_333
timestamp 0
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_345
timestamp 0
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_357
timestamp 0
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_363
timestamp 0
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_365
timestamp 0
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_377
timestamp 0
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_389
timestamp 0
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_401
timestamp 0
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_413
timestamp 0
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_419
timestamp 0
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_421
timestamp 0
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_433
timestamp 0
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_445
timestamp 0
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_457
timestamp 0
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_469
timestamp 0
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_475
timestamp 0
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_477
timestamp 0
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_489
timestamp 0
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_501
timestamp 0
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_513
timestamp 0
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_525
timestamp 0
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_531
timestamp 0
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_533
timestamp 0
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_545
timestamp 0
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_557
timestamp 0
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_569
timestamp 0
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_581
timestamp 0
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_587
timestamp 0
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_589
timestamp 0
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_601
timestamp 0
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_613
timestamp 0
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_3
timestamp 0
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_15
timestamp 0
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_27
timestamp 0
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_39
timestamp 0
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_51
timestamp 0
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_55
timestamp 0
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_57
timestamp 0
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_69
timestamp 0
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_81
timestamp 0
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_93
timestamp 0
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_105
timestamp 0
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_111
timestamp 0
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_113
timestamp 0
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_125
timestamp 0
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_137
timestamp 0
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_149
timestamp 0
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_161
timestamp 0
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_167
timestamp 0
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_169
timestamp 0
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_181
timestamp 0
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_193
timestamp 0
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_205
timestamp 0
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_217
timestamp 0
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_223
timestamp 0
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_225
timestamp 0
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_237
timestamp 0
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_249
timestamp 0
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_261
timestamp 0
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_273
timestamp 0
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_279
timestamp 0
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_281
timestamp 0
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_293
timestamp 0
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_305
timestamp 0
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_317
timestamp 0
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_329
timestamp 0
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_335
timestamp 0
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_337
timestamp 0
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_349
timestamp 0
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_361
timestamp 0
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_373
timestamp 0
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_385
timestamp 0
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_391
timestamp 0
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_393
timestamp 0
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_405
timestamp 0
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_417
timestamp 0
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_429
timestamp 0
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_441
timestamp 0
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_447
timestamp 0
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_449
timestamp 0
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_461
timestamp 0
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_473
timestamp 0
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_485
timestamp 0
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_497
timestamp 0
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_503
timestamp 0
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_505
timestamp 0
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_517
timestamp 0
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_529
timestamp 0
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_541
timestamp 0
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_553
timestamp 0
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_559
timestamp 0
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_561
timestamp 0
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_573
timestamp 0
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_585
timestamp 0
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_597
timestamp 0
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_609
timestamp 0
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_615
timestamp 0
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_617
timestamp 0
transform 1 0 57868 0 -1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_3
timestamp 0
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_15
timestamp 0
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_27
timestamp 0
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_29
timestamp 0
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_41
timestamp 0
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_53
timestamp 0
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_65
timestamp 0
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_77
timestamp 0
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_83
timestamp 0
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_85
timestamp 0
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_97
timestamp 0
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_109
timestamp 0
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_121
timestamp 0
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_133
timestamp 0
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_139
timestamp 0
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_141
timestamp 0
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_153
timestamp 0
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_165
timestamp 0
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_177
timestamp 0
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_189
timestamp 0
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_195
timestamp 0
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_197
timestamp 0
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_209
timestamp 0
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_221
timestamp 0
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_233
timestamp 0
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_245
timestamp 0
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_251
timestamp 0
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_253
timestamp 0
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_265
timestamp 0
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_277
timestamp 0
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_289
timestamp 0
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_301
timestamp 0
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_307
timestamp 0
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_309
timestamp 0
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_321
timestamp 0
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_333
timestamp 0
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_345
timestamp 0
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_357
timestamp 0
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_363
timestamp 0
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_365
timestamp 0
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_377
timestamp 0
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_389
timestamp 0
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_401
timestamp 0
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_413
timestamp 0
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_419
timestamp 0
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_421
timestamp 0
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_433
timestamp 0
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_445
timestamp 0
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_457
timestamp 0
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_469
timestamp 0
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_475
timestamp 0
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_477
timestamp 0
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_489
timestamp 0
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_501
timestamp 0
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_513
timestamp 0
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_525
timestamp 0
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_531
timestamp 0
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_533
timestamp 0
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_545
timestamp 0
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_557
timestamp 0
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_569
timestamp 0
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_581
timestamp 0
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_587
timestamp 0
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_589
timestamp 0
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_601
timestamp 0
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_613
timestamp 0
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_3
timestamp 0
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_15
timestamp 0
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_27
timestamp 0
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_39
timestamp 0
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_51
timestamp 0
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_55
timestamp 0
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_57
timestamp 0
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_69
timestamp 0
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_81
timestamp 0
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_93
timestamp 0
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_105
timestamp 0
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_111
timestamp 0
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_113
timestamp 0
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_125
timestamp 0
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_137
timestamp 0
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_149
timestamp 0
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_161
timestamp 0
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_167
timestamp 0
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_169
timestamp 0
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_181
timestamp 0
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_193
timestamp 0
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_205
timestamp 0
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_217
timestamp 0
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_223
timestamp 0
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_225
timestamp 0
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_237
timestamp 0
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_249
timestamp 0
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_261
timestamp 0
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_273
timestamp 0
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_279
timestamp 0
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_281
timestamp 0
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_293
timestamp 0
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_305
timestamp 0
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_317
timestamp 0
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_329
timestamp 0
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_335
timestamp 0
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_337
timestamp 0
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_349
timestamp 0
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_361
timestamp 0
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_373
timestamp 0
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_385
timestamp 0
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_391
timestamp 0
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_393
timestamp 0
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_405
timestamp 0
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_417
timestamp 0
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_429
timestamp 0
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_441
timestamp 0
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_447
timestamp 0
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_449
timestamp 0
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_461
timestamp 0
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_473
timestamp 0
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_485
timestamp 0
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_497
timestamp 0
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_503
timestamp 0
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_505
timestamp 0
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_517
timestamp 0
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_529
timestamp 0
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_541
timestamp 0
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_553
timestamp 0
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_559
timestamp 0
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_561
timestamp 0
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_573
timestamp 0
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_585
timestamp 0
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_597
timestamp 0
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_609
timestamp 0
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_615
timestamp 0
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_617
timestamp 0
transform 1 0 57868 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_3
timestamp 0
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_15
timestamp 0
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_27
timestamp 0
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_29
timestamp 0
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_41
timestamp 0
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_53
timestamp 0
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_65
timestamp 0
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_77
timestamp 0
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_83
timestamp 0
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_85
timestamp 0
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_97
timestamp 0
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_109
timestamp 0
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_121
timestamp 0
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_133
timestamp 0
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_139
timestamp 0
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_141
timestamp 0
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_153
timestamp 0
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_165
timestamp 0
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_177
timestamp 0
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_189
timestamp 0
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_195
timestamp 0
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_197
timestamp 0
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_209
timestamp 0
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_221
timestamp 0
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_233
timestamp 0
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_245
timestamp 0
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_251
timestamp 0
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_253
timestamp 0
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_265
timestamp 0
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_277
timestamp 0
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_289
timestamp 0
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_301
timestamp 0
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_307
timestamp 0
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_309
timestamp 0
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_321
timestamp 0
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_333
timestamp 0
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_345
timestamp 0
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_357
timestamp 0
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_363
timestamp 0
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_365
timestamp 0
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_377
timestamp 0
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_389
timestamp 0
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_401
timestamp 0
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_413
timestamp 0
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_419
timestamp 0
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_421
timestamp 0
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_433
timestamp 0
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_445
timestamp 0
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_457
timestamp 0
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_469
timestamp 0
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_475
timestamp 0
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_477
timestamp 0
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_489
timestamp 0
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_501
timestamp 0
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_513
timestamp 0
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_525
timestamp 0
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_531
timestamp 0
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_533
timestamp 0
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_545
timestamp 0
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_557
timestamp 0
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_569
timestamp 0
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_581
timestamp 0
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_587
timestamp 0
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_589
timestamp 0
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_601
timestamp 0
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_613
timestamp 0
transform 1 0 57500 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_3
timestamp 0
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_15
timestamp 0
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_27
timestamp 0
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_39
timestamp 0
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_51
timestamp 0
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_55
timestamp 0
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_57
timestamp 0
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_69
timestamp 0
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_81
timestamp 0
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_93
timestamp 0
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_105
timestamp 0
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_111
timestamp 0
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_113
timestamp 0
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_125
timestamp 0
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_137
timestamp 0
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_149
timestamp 0
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_161
timestamp 0
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_167
timestamp 0
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_169
timestamp 0
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_181
timestamp 0
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_193
timestamp 0
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_205
timestamp 0
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_217
timestamp 0
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_223
timestamp 0
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_225
timestamp 0
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_237
timestamp 0
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_249
timestamp 0
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_261
timestamp 0
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_273
timestamp 0
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_279
timestamp 0
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_281
timestamp 0
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_293
timestamp 0
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_305
timestamp 0
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_317
timestamp 0
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_329
timestamp 0
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_335
timestamp 0
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_337
timestamp 0
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_349
timestamp 0
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_361
timestamp 0
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_373
timestamp 0
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_385
timestamp 0
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_391
timestamp 0
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_393
timestamp 0
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_405
timestamp 0
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_417
timestamp 0
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_429
timestamp 0
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_441
timestamp 0
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_447
timestamp 0
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_449
timestamp 0
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_461
timestamp 0
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_473
timestamp 0
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_485
timestamp 0
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_497
timestamp 0
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_503
timestamp 0
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_505
timestamp 0
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_517
timestamp 0
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_529
timestamp 0
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_541
timestamp 0
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_553
timestamp 0
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_559
timestamp 0
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_561
timestamp 0
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_573
timestamp 0
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_585
timestamp 0
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_597
timestamp 0
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_609
timestamp 0
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_615
timestamp 0
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_617
timestamp 0
transform 1 0 57868 0 -1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_3
timestamp 0
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_15
timestamp 0
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_27
timestamp 0
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_29
timestamp 0
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_41
timestamp 0
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_53
timestamp 0
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_65
timestamp 0
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_77
timestamp 0
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_83
timestamp 0
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_85
timestamp 0
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_97
timestamp 0
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_109
timestamp 0
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_121
timestamp 0
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_133
timestamp 0
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_139
timestamp 0
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_141
timestamp 0
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_153
timestamp 0
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_165
timestamp 0
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_177
timestamp 0
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_189
timestamp 0
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_195
timestamp 0
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_197
timestamp 0
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_209
timestamp 0
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_221
timestamp 0
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_233
timestamp 0
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_245
timestamp 0
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_251
timestamp 0
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_253
timestamp 0
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_265
timestamp 0
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_277
timestamp 0
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_289
timestamp 0
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_301
timestamp 0
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_307
timestamp 0
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_309
timestamp 0
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_321
timestamp 0
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_333
timestamp 0
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_345
timestamp 0
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_357
timestamp 0
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_363
timestamp 0
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_365
timestamp 0
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_377
timestamp 0
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_389
timestamp 0
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_401
timestamp 0
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_413
timestamp 0
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_419
timestamp 0
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_421
timestamp 0
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_433
timestamp 0
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_445
timestamp 0
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_457
timestamp 0
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_469
timestamp 0
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_475
timestamp 0
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_477
timestamp 0
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_489
timestamp 0
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_501
timestamp 0
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_513
timestamp 0
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_525
timestamp 0
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_531
timestamp 0
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_533
timestamp 0
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_545
timestamp 0
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_557
timestamp 0
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_569
timestamp 0
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_581
timestamp 0
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_587
timestamp 0
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_589
timestamp 0
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_601
timestamp 0
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_613
timestamp 0
transform 1 0 57500 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_3
timestamp 0
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_15
timestamp 0
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_27
timestamp 0
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_39
timestamp 0
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_51
timestamp 0
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_55
timestamp 0
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_57
timestamp 0
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_69
timestamp 0
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_81
timestamp 0
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_93
timestamp 0
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_105
timestamp 0
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_111
timestamp 0
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_113
timestamp 0
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_125
timestamp 0
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_137
timestamp 0
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_149
timestamp 0
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_161
timestamp 0
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_167
timestamp 0
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_169
timestamp 0
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_181
timestamp 0
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_193
timestamp 0
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_205
timestamp 0
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_217
timestamp 0
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_223
timestamp 0
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_225
timestamp 0
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_237
timestamp 0
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_249
timestamp 0
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_261
timestamp 0
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_273
timestamp 0
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_279
timestamp 0
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_281
timestamp 0
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_293
timestamp 0
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_305
timestamp 0
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_317
timestamp 0
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_329
timestamp 0
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_335
timestamp 0
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_337
timestamp 0
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_349
timestamp 0
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_361
timestamp 0
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_373
timestamp 0
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_385
timestamp 0
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_391
timestamp 0
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_393
timestamp 0
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_405
timestamp 0
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_417
timestamp 0
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_429
timestamp 0
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_441
timestamp 0
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_447
timestamp 0
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_449
timestamp 0
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_461
timestamp 0
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_473
timestamp 0
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_485
timestamp 0
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_497
timestamp 0
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_503
timestamp 0
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_505
timestamp 0
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_517
timestamp 0
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_529
timestamp 0
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_541
timestamp 0
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_553
timestamp 0
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_559
timestamp 0
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_561
timestamp 0
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_573
timestamp 0
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_585
timestamp 0
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_597
timestamp 0
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_609
timestamp 0
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_615
timestamp 0
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_617
timestamp 0
transform 1 0 57868 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_3
timestamp 0
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_15
timestamp 0
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_27
timestamp 0
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_29
timestamp 0
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_41
timestamp 0
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_53
timestamp 0
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_65
timestamp 0
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_77
timestamp 0
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_83
timestamp 0
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_85
timestamp 0
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_97
timestamp 0
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_109
timestamp 0
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_121
timestamp 0
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_133
timestamp 0
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_139
timestamp 0
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_141
timestamp 0
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_153
timestamp 0
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_165
timestamp 0
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_177
timestamp 0
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_189
timestamp 0
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_195
timestamp 0
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_197
timestamp 0
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_209
timestamp 0
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_221
timestamp 0
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_233
timestamp 0
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_245
timestamp 0
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_251
timestamp 0
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_253
timestamp 0
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_265
timestamp 0
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_277
timestamp 0
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_289
timestamp 0
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_301
timestamp 0
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_307
timestamp 0
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_309
timestamp 0
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_321
timestamp 0
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_333
timestamp 0
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_345
timestamp 0
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_357
timestamp 0
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_363
timestamp 0
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_365
timestamp 0
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_377
timestamp 0
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_389
timestamp 0
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_401
timestamp 0
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_413
timestamp 0
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_419
timestamp 0
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_421
timestamp 0
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_433
timestamp 0
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_445
timestamp 0
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_457
timestamp 0
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_469
timestamp 0
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_475
timestamp 0
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_477
timestamp 0
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_489
timestamp 0
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_501
timestamp 0
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_513
timestamp 0
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_525
timestamp 0
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_531
timestamp 0
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_533
timestamp 0
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_545
timestamp 0
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_557
timestamp 0
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_569
timestamp 0
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_581
timestamp 0
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_587
timestamp 0
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_589
timestamp 0
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_601
timestamp 0
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_613
timestamp 0
transform 1 0 57500 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_3
timestamp 0
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_15
timestamp 0
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_27
timestamp 0
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_39
timestamp 0
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_51
timestamp 0
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_55
timestamp 0
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_57
timestamp 0
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_69
timestamp 0
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_81
timestamp 0
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_93
timestamp 0
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_105
timestamp 0
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_111
timestamp 0
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_113
timestamp 0
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_125
timestamp 0
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_137
timestamp 0
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_149
timestamp 0
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_161
timestamp 0
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_167
timestamp 0
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_169
timestamp 0
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_181
timestamp 0
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_193
timestamp 0
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_205
timestamp 0
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_217
timestamp 0
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_223
timestamp 0
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_225
timestamp 0
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_237
timestamp 0
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_249
timestamp 0
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_261
timestamp 0
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_273
timestamp 0
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_279
timestamp 0
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_281
timestamp 0
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_293
timestamp 0
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_305
timestamp 0
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_317
timestamp 0
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_329
timestamp 0
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_335
timestamp 0
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_337
timestamp 0
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_349
timestamp 0
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_361
timestamp 0
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_373
timestamp 0
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_385
timestamp 0
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_391
timestamp 0
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_393
timestamp 0
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_405
timestamp 0
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_417
timestamp 0
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_429
timestamp 0
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_441
timestamp 0
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_447
timestamp 0
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_449
timestamp 0
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_461
timestamp 0
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_473
timestamp 0
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_485
timestamp 0
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_497
timestamp 0
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_503
timestamp 0
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_505
timestamp 0
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_517
timestamp 0
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_529
timestamp 0
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_541
timestamp 0
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_553
timestamp 0
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_559
timestamp 0
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_561
timestamp 0
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_573
timestamp 0
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_585
timestamp 0
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_597
timestamp 0
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_609
timestamp 0
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_615
timestamp 0
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_617
timestamp 0
transform 1 0 57868 0 -1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_3
timestamp 0
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_15
timestamp 0
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_27
timestamp 0
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_29
timestamp 0
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_41
timestamp 0
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_53
timestamp 0
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_65
timestamp 0
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_77
timestamp 0
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_83
timestamp 0
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_85
timestamp 0
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_97
timestamp 0
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_109
timestamp 0
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_121
timestamp 0
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_133
timestamp 0
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_139
timestamp 0
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_141
timestamp 0
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_153
timestamp 0
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_165
timestamp 0
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_177
timestamp 0
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_189
timestamp 0
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_195
timestamp 0
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_197
timestamp 0
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_209
timestamp 0
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_221
timestamp 0
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_233
timestamp 0
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_245
timestamp 0
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_251
timestamp 0
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_253
timestamp 0
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_265
timestamp 0
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_277
timestamp 0
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_289
timestamp 0
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_301
timestamp 0
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_307
timestamp 0
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_309
timestamp 0
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_321
timestamp 0
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_333
timestamp 0
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_345
timestamp 0
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_357
timestamp 0
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_363
timestamp 0
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_365
timestamp 0
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_377
timestamp 0
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_389
timestamp 0
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_401
timestamp 0
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_413
timestamp 0
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_419
timestamp 0
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_421
timestamp 0
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_433
timestamp 0
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_445
timestamp 0
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_457
timestamp 0
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_469
timestamp 0
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_475
timestamp 0
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_477
timestamp 0
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_489
timestamp 0
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_501
timestamp 0
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_513
timestamp 0
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_525
timestamp 0
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_531
timestamp 0
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_533
timestamp 0
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_545
timestamp 0
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_557
timestamp 0
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_569
timestamp 0
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_581
timestamp 0
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_587
timestamp 0
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_589
timestamp 0
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_601
timestamp 0
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_613
timestamp 0
transform 1 0 57500 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_3
timestamp 0
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_15
timestamp 0
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_27
timestamp 0
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_39
timestamp 0
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_51
timestamp 0
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_55
timestamp 0
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_57
timestamp 0
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_69
timestamp 0
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_81
timestamp 0
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_93
timestamp 0
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_105
timestamp 0
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_111
timestamp 0
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_113
timestamp 0
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_125
timestamp 0
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_137
timestamp 0
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_149
timestamp 0
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_161
timestamp 0
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_167
timestamp 0
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_169
timestamp 0
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_181
timestamp 0
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_193
timestamp 0
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_205
timestamp 0
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_217
timestamp 0
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_223
timestamp 0
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_225
timestamp 0
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_237
timestamp 0
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_249
timestamp 0
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_261
timestamp 0
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_273
timestamp 0
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_279
timestamp 0
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_281
timestamp 0
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_293
timestamp 0
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_305
timestamp 0
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_317
timestamp 0
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_329
timestamp 0
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_335
timestamp 0
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_337
timestamp 0
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_349
timestamp 0
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_361
timestamp 0
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_373
timestamp 0
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_385
timestamp 0
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_391
timestamp 0
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_393
timestamp 0
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_405
timestamp 0
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_417
timestamp 0
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_429
timestamp 0
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_441
timestamp 0
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_447
timestamp 0
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_449
timestamp 0
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_461
timestamp 0
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_473
timestamp 0
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_485
timestamp 0
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_497
timestamp 0
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_503
timestamp 0
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_505
timestamp 0
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_517
timestamp 0
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_529
timestamp 0
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_541
timestamp 0
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_553
timestamp 0
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_559
timestamp 0
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_561
timestamp 0
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_573
timestamp 0
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_585
timestamp 0
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_597
timestamp 0
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_609
timestamp 0
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_615
timestamp 0
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_617
timestamp 0
transform 1 0 57868 0 -1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_3
timestamp 0
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_15
timestamp 0
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_27
timestamp 0
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_29
timestamp 0
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_41
timestamp 0
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_53
timestamp 0
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_65
timestamp 0
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_77
timestamp 0
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_83
timestamp 0
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_85
timestamp 0
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_97
timestamp 0
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_109
timestamp 0
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_121
timestamp 0
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_133
timestamp 0
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_139
timestamp 0
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_141
timestamp 0
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_153
timestamp 0
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_165
timestamp 0
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_177
timestamp 0
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_189
timestamp 0
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_195
timestamp 0
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_197
timestamp 0
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_209
timestamp 0
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_221
timestamp 0
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_233
timestamp 0
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_245
timestamp 0
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_251
timestamp 0
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_253
timestamp 0
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_265
timestamp 0
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_277
timestamp 0
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_289
timestamp 0
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_301
timestamp 0
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_307
timestamp 0
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_309
timestamp 0
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_321
timestamp 0
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_333
timestamp 0
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_345
timestamp 0
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_357
timestamp 0
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_363
timestamp 0
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_365
timestamp 0
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_377
timestamp 0
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_389
timestamp 0
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_401
timestamp 0
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_413
timestamp 0
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_419
timestamp 0
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_421
timestamp 0
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_433
timestamp 0
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_445
timestamp 0
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_457
timestamp 0
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_469
timestamp 0
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_475
timestamp 0
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_477
timestamp 0
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_489
timestamp 0
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_501
timestamp 0
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_513
timestamp 0
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_525
timestamp 0
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_531
timestamp 0
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_533
timestamp 0
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_545
timestamp 0
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_557
timestamp 0
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_569
timestamp 0
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_581
timestamp 0
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_587
timestamp 0
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_589
timestamp 0
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_601
timestamp 0
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_613
timestamp 0
transform 1 0 57500 0 1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_3
timestamp 0
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_15
timestamp 0
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_27
timestamp 0
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_39
timestamp 0
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_51
timestamp 0
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_55
timestamp 0
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_57
timestamp 0
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_69
timestamp 0
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_81
timestamp 0
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_93
timestamp 0
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_105
timestamp 0
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_111
timestamp 0
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_113
timestamp 0
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_125
timestamp 0
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_137
timestamp 0
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_149
timestamp 0
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_161
timestamp 0
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_167
timestamp 0
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_169
timestamp 0
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_181
timestamp 0
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_193
timestamp 0
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_205
timestamp 0
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_217
timestamp 0
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_223
timestamp 0
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_225
timestamp 0
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_237
timestamp 0
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_249
timestamp 0
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_261
timestamp 0
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_273
timestamp 0
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_279
timestamp 0
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_281
timestamp 0
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_293
timestamp 0
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_305
timestamp 0
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_317
timestamp 0
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_329
timestamp 0
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_335
timestamp 0
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_337
timestamp 0
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_349
timestamp 0
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_361
timestamp 0
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_373
timestamp 0
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_385
timestamp 0
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_391
timestamp 0
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_393
timestamp 0
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_405
timestamp 0
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_417
timestamp 0
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_429
timestamp 0
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_441
timestamp 0
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_447
timestamp 0
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_449
timestamp 0
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_461
timestamp 0
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_473
timestamp 0
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_485
timestamp 0
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_497
timestamp 0
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_503
timestamp 0
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_505
timestamp 0
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_517
timestamp 0
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_529
timestamp 0
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_541
timestamp 0
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_553
timestamp 0
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_559
timestamp 0
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_561
timestamp 0
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_573
timestamp 0
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_585
timestamp 0
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_597
timestamp 0
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_609
timestamp 0
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_615
timestamp 0
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_617
timestamp 0
transform 1 0 57868 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_3
timestamp 0
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_15
timestamp 0
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_27
timestamp 0
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_29
timestamp 0
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_41
timestamp 0
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_53
timestamp 0
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_65
timestamp 0
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_77
timestamp 0
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_83
timestamp 0
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_85
timestamp 0
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_97
timestamp 0
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_109
timestamp 0
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_121
timestamp 0
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_133
timestamp 0
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_139
timestamp 0
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_141
timestamp 0
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_153
timestamp 0
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_165
timestamp 0
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_177
timestamp 0
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_189
timestamp 0
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_195
timestamp 0
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_197
timestamp 0
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_209
timestamp 0
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_221
timestamp 0
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_233
timestamp 0
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_245
timestamp 0
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_251
timestamp 0
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_253
timestamp 0
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_265
timestamp 0
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_277
timestamp 0
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_289
timestamp 0
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_301
timestamp 0
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_307
timestamp 0
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_309
timestamp 0
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_321
timestamp 0
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_333
timestamp 0
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_345
timestamp 0
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_357
timestamp 0
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_363
timestamp 0
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_365
timestamp 0
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_377
timestamp 0
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_389
timestamp 0
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_401
timestamp 0
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_413
timestamp 0
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_419
timestamp 0
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_421
timestamp 0
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_433
timestamp 0
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_445
timestamp 0
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_457
timestamp 0
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_469
timestamp 0
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_475
timestamp 0
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_477
timestamp 0
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_489
timestamp 0
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_501
timestamp 0
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_513
timestamp 0
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_525
timestamp 0
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_531
timestamp 0
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_533
timestamp 0
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_545
timestamp 0
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_557
timestamp 0
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_569
timestamp 0
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_581
timestamp 0
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_587
timestamp 0
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_589
timestamp 0
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_601
timestamp 0
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_613
timestamp 0
transform 1 0 57500 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_3
timestamp 0
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_15
timestamp 0
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_27
timestamp 0
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_39
timestamp 0
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_81_51
timestamp 0
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_55
timestamp 0
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_57
timestamp 0
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_69
timestamp 0
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_81
timestamp 0
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_93
timestamp 0
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_105
timestamp 0
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_111
timestamp 0
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_113
timestamp 0
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_125
timestamp 0
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_137
timestamp 0
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_149
timestamp 0
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_161
timestamp 0
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_167
timestamp 0
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_169
timestamp 0
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_181
timestamp 0
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_193
timestamp 0
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_205
timestamp 0
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_217
timestamp 0
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_223
timestamp 0
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_225
timestamp 0
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_237
timestamp 0
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_249
timestamp 0
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_261
timestamp 0
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_273
timestamp 0
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_279
timestamp 0
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_281
timestamp 0
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_293
timestamp 0
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_305
timestamp 0
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_317
timestamp 0
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_329
timestamp 0
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_335
timestamp 0
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_337
timestamp 0
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_349
timestamp 0
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_361
timestamp 0
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_373
timestamp 0
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_385
timestamp 0
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_391
timestamp 0
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_393
timestamp 0
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_405
timestamp 0
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_417
timestamp 0
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_429
timestamp 0
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_441
timestamp 0
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_447
timestamp 0
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_449
timestamp 0
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_461
timestamp 0
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_473
timestamp 0
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_485
timestamp 0
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_497
timestamp 0
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_503
timestamp 0
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_505
timestamp 0
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_517
timestamp 0
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_529
timestamp 0
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_541
timestamp 0
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_553
timestamp 0
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_559
timestamp 0
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_561
timestamp 0
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_573
timestamp 0
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_585
timestamp 0
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_597
timestamp 0
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_609
timestamp 0
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_615
timestamp 0
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_81_617
timestamp 0
transform 1 0 57868 0 -1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_3
timestamp 0
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_15
timestamp 0
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_27
timestamp 0
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_29
timestamp 0
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_41
timestamp 0
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_53
timestamp 0
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_65
timestamp 0
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_77
timestamp 0
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_83
timestamp 0
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_85
timestamp 0
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_97
timestamp 0
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_109
timestamp 0
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_121
timestamp 0
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_133
timestamp 0
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_139
timestamp 0
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_141
timestamp 0
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_153
timestamp 0
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_165
timestamp 0
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_177
timestamp 0
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_189
timestamp 0
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_195
timestamp 0
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_197
timestamp 0
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_209
timestamp 0
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_221
timestamp 0
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_233
timestamp 0
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_245
timestamp 0
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_251
timestamp 0
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_253
timestamp 0
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_265
timestamp 0
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_277
timestamp 0
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_289
timestamp 0
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_301
timestamp 0
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_307
timestamp 0
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_309
timestamp 0
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_321
timestamp 0
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_333
timestamp 0
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_345
timestamp 0
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_357
timestamp 0
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_363
timestamp 0
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_365
timestamp 0
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_377
timestamp 0
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_389
timestamp 0
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_401
timestamp 0
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_413
timestamp 0
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_419
timestamp 0
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_421
timestamp 0
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_433
timestamp 0
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_445
timestamp 0
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_457
timestamp 0
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_469
timestamp 0
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_475
timestamp 0
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_477
timestamp 0
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_489
timestamp 0
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_501
timestamp 0
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_513
timestamp 0
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_525
timestamp 0
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_531
timestamp 0
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_533
timestamp 0
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_545
timestamp 0
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_557
timestamp 0
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_569
timestamp 0
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_581
timestamp 0
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_587
timestamp 0
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_589
timestamp 0
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_601
timestamp 0
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_613
timestamp 0
transform 1 0 57500 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_3
timestamp 0
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_15
timestamp 0
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_27
timestamp 0
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_39
timestamp 0
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83_51
timestamp 0
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_55
timestamp 0
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_57
timestamp 0
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_69
timestamp 0
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_81
timestamp 0
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_93
timestamp 0
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_105
timestamp 0
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_111
timestamp 0
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_113
timestamp 0
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_125
timestamp 0
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_137
timestamp 0
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_149
timestamp 0
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_161
timestamp 0
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_167
timestamp 0
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_169
timestamp 0
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_181
timestamp 0
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_193
timestamp 0
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_205
timestamp 0
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_217
timestamp 0
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_223
timestamp 0
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_225
timestamp 0
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_237
timestamp 0
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_249
timestamp 0
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_261
timestamp 0
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_273
timestamp 0
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_279
timestamp 0
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_281
timestamp 0
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_293
timestamp 0
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_305
timestamp 0
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_317
timestamp 0
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_329
timestamp 0
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_335
timestamp 0
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_337
timestamp 0
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_349
timestamp 0
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_361
timestamp 0
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_373
timestamp 0
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_385
timestamp 0
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_391
timestamp 0
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_393
timestamp 0
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_405
timestamp 0
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_417
timestamp 0
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_429
timestamp 0
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_441
timestamp 0
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_447
timestamp 0
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_449
timestamp 0
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_461
timestamp 0
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_473
timestamp 0
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_485
timestamp 0
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_497
timestamp 0
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_503
timestamp 0
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_505
timestamp 0
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_517
timestamp 0
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_529
timestamp 0
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_541
timestamp 0
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_553
timestamp 0
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_559
timestamp 0
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_561
timestamp 0
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_573
timestamp 0
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_585
timestamp 0
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_597
timestamp 0
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_609
timestamp 0
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_615
timestamp 0
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_83_617
timestamp 0
transform 1 0 57868 0 -1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_3
timestamp 0
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_15
timestamp 0
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_27
timestamp 0
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_29
timestamp 0
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_41
timestamp 0
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_53
timestamp 0
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_65
timestamp 0
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_77
timestamp 0
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_83
timestamp 0
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_85
timestamp 0
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_97
timestamp 0
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_109
timestamp 0
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_121
timestamp 0
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_133
timestamp 0
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_139
timestamp 0
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_141
timestamp 0
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_153
timestamp 0
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_165
timestamp 0
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_177
timestamp 0
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_189
timestamp 0
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_195
timestamp 0
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_197
timestamp 0
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_209
timestamp 0
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_221
timestamp 0
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_233
timestamp 0
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_245
timestamp 0
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_251
timestamp 0
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_253
timestamp 0
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_265
timestamp 0
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_277
timestamp 0
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_289
timestamp 0
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_301
timestamp 0
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_307
timestamp 0
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_309
timestamp 0
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_321
timestamp 0
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_333
timestamp 0
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_345
timestamp 0
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_357
timestamp 0
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_363
timestamp 0
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_365
timestamp 0
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_377
timestamp 0
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_389
timestamp 0
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_401
timestamp 0
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_413
timestamp 0
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_419
timestamp 0
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_421
timestamp 0
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_433
timestamp 0
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_445
timestamp 0
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_457
timestamp 0
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_469
timestamp 0
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_475
timestamp 0
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_477
timestamp 0
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_489
timestamp 0
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_501
timestamp 0
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_513
timestamp 0
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_525
timestamp 0
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_531
timestamp 0
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_533
timestamp 0
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_545
timestamp 0
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_557
timestamp 0
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_569
timestamp 0
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_581
timestamp 0
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_587
timestamp 0
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_589
timestamp 0
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_601
timestamp 0
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_613
timestamp 0
transform 1 0 57500 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_3
timestamp 0
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_15
timestamp 0
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_27
timestamp 0
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_39
timestamp 0
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85_51
timestamp 0
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_55
timestamp 0
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_57
timestamp 0
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_69
timestamp 0
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_81
timestamp 0
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_93
timestamp 0
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_105
timestamp 0
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_111
timestamp 0
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_113
timestamp 0
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_125
timestamp 0
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_137
timestamp 0
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_149
timestamp 0
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_161
timestamp 0
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_167
timestamp 0
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_169
timestamp 0
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_181
timestamp 0
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_193
timestamp 0
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_205
timestamp 0
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_217
timestamp 0
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_223
timestamp 0
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_225
timestamp 0
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_237
timestamp 0
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_249
timestamp 0
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_261
timestamp 0
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_273
timestamp 0
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_279
timestamp 0
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_281
timestamp 0
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_293
timestamp 0
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_305
timestamp 0
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_317
timestamp 0
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_329
timestamp 0
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_335
timestamp 0
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_337
timestamp 0
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_349
timestamp 0
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_361
timestamp 0
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_373
timestamp 0
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_385
timestamp 0
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_391
timestamp 0
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_393
timestamp 0
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_405
timestamp 0
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_417
timestamp 0
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_429
timestamp 0
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_441
timestamp 0
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_447
timestamp 0
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_449
timestamp 0
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_461
timestamp 0
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_473
timestamp 0
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_485
timestamp 0
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_497
timestamp 0
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_503
timestamp 0
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_505
timestamp 0
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_517
timestamp 0
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_529
timestamp 0
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_541
timestamp 0
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_553
timestamp 0
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_559
timestamp 0
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_561
timestamp 0
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_573
timestamp 0
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_585
timestamp 0
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_597
timestamp 0
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_609
timestamp 0
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_615
timestamp 0
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85_617
timestamp 0
transform 1 0 57868 0 -1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_3
timestamp 0
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_15
timestamp 0
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_27
timestamp 0
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_29
timestamp 0
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_41
timestamp 0
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_53
timestamp 0
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_65
timestamp 0
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_77
timestamp 0
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_83
timestamp 0
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_85
timestamp 0
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_97
timestamp 0
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_109
timestamp 0
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_121
timestamp 0
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_133
timestamp 0
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_139
timestamp 0
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_141
timestamp 0
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_153
timestamp 0
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_165
timestamp 0
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_177
timestamp 0
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_189
timestamp 0
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_195
timestamp 0
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_197
timestamp 0
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_209
timestamp 0
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_221
timestamp 0
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_233
timestamp 0
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_245
timestamp 0
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_251
timestamp 0
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_253
timestamp 0
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_265
timestamp 0
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_277
timestamp 0
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_289
timestamp 0
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_301
timestamp 0
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_307
timestamp 0
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_309
timestamp 0
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_321
timestamp 0
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_333
timestamp 0
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_345
timestamp 0
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_357
timestamp 0
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_363
timestamp 0
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_365
timestamp 0
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_377
timestamp 0
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_389
timestamp 0
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_401
timestamp 0
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_413
timestamp 0
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_419
timestamp 0
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_421
timestamp 0
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_433
timestamp 0
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_445
timestamp 0
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_457
timestamp 0
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_469
timestamp 0
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_475
timestamp 0
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_477
timestamp 0
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_489
timestamp 0
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_501
timestamp 0
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_513
timestamp 0
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_525
timestamp 0
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_531
timestamp 0
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_533
timestamp 0
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_545
timestamp 0
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_557
timestamp 0
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_569
timestamp 0
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_581
timestamp 0
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_587
timestamp 0
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_589
timestamp 0
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_601
timestamp 0
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_613
timestamp 0
transform 1 0 57500 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_3
timestamp 0
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_15
timestamp 0
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_27
timestamp 0
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_39
timestamp 0
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_87_51
timestamp 0
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_55
timestamp 0
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_57
timestamp 0
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_69
timestamp 0
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_81
timestamp 0
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_93
timestamp 0
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_105
timestamp 0
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_111
timestamp 0
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_113
timestamp 0
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_125
timestamp 0
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_137
timestamp 0
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_149
timestamp 0
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_161
timestamp 0
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_167
timestamp 0
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_169
timestamp 0
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_181
timestamp 0
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_193
timestamp 0
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_205
timestamp 0
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_217
timestamp 0
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_223
timestamp 0
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_225
timestamp 0
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_237
timestamp 0
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_249
timestamp 0
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_261
timestamp 0
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_273
timestamp 0
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_279
timestamp 0
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_281
timestamp 0
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_293
timestamp 0
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_305
timestamp 0
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_317
timestamp 0
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_329
timestamp 0
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_335
timestamp 0
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_337
timestamp 0
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_349
timestamp 0
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_361
timestamp 0
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_373
timestamp 0
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_385
timestamp 0
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_391
timestamp 0
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_393
timestamp 0
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_405
timestamp 0
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_417
timestamp 0
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_429
timestamp 0
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_441
timestamp 0
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_447
timestamp 0
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_449
timestamp 0
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_461
timestamp 0
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_473
timestamp 0
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_485
timestamp 0
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_497
timestamp 0
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_503
timestamp 0
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_505
timestamp 0
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_517
timestamp 0
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_529
timestamp 0
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_541
timestamp 0
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_553
timestamp 0
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_559
timestamp 0
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_561
timestamp 0
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_573
timestamp 0
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_585
timestamp 0
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_597
timestamp 0
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_609
timestamp 0
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_615
timestamp 0
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_87_617
timestamp 0
transform 1 0 57868 0 -1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_3
timestamp 0
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_15
timestamp 0
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_27
timestamp 0
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_29
timestamp 0
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_41
timestamp 0
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_53
timestamp 0
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_65
timestamp 0
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_77
timestamp 0
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_83
timestamp 0
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_85
timestamp 0
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_97
timestamp 0
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_109
timestamp 0
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_121
timestamp 0
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_133
timestamp 0
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_139
timestamp 0
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_141
timestamp 0
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_153
timestamp 0
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_165
timestamp 0
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_177
timestamp 0
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_189
timestamp 0
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_195
timestamp 0
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_197
timestamp 0
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_209
timestamp 0
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_221
timestamp 0
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_233
timestamp 0
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_245
timestamp 0
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_251
timestamp 0
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_253
timestamp 0
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_265
timestamp 0
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_277
timestamp 0
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_289
timestamp 0
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_301
timestamp 0
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_307
timestamp 0
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_309
timestamp 0
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_321
timestamp 0
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_333
timestamp 0
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_345
timestamp 0
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_357
timestamp 0
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_363
timestamp 0
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_365
timestamp 0
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_377
timestamp 0
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_389
timestamp 0
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_401
timestamp 0
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_413
timestamp 0
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_419
timestamp 0
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_421
timestamp 0
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_433
timestamp 0
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_445
timestamp 0
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_457
timestamp 0
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_469
timestamp 0
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_475
timestamp 0
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_477
timestamp 0
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_489
timestamp 0
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_501
timestamp 0
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_513
timestamp 0
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_525
timestamp 0
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_531
timestamp 0
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_533
timestamp 0
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_545
timestamp 0
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_557
timestamp 0
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_569
timestamp 0
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_581
timestamp 0
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_587
timestamp 0
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_589
timestamp 0
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_601
timestamp 0
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_613
timestamp 0
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_3
timestamp 0
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_15
timestamp 0
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_27
timestamp 0
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_39
timestamp 0
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89_51
timestamp 0
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_55
timestamp 0
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_57
timestamp 0
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_69
timestamp 0
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_81
timestamp 0
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_93
timestamp 0
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_105
timestamp 0
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_111
timestamp 0
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_113
timestamp 0
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_125
timestamp 0
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_137
timestamp 0
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_149
timestamp 0
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_161
timestamp 0
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_167
timestamp 0
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_169
timestamp 0
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_181
timestamp 0
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_193
timestamp 0
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_205
timestamp 0
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_217
timestamp 0
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_223
timestamp 0
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_225
timestamp 0
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_237
timestamp 0
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_249
timestamp 0
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_261
timestamp 0
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_273
timestamp 0
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_279
timestamp 0
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_281
timestamp 0
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_293
timestamp 0
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_305
timestamp 0
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_317
timestamp 0
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_329
timestamp 0
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_335
timestamp 0
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_337
timestamp 0
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_349
timestamp 0
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_361
timestamp 0
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_373
timestamp 0
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_385
timestamp 0
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_391
timestamp 0
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_393
timestamp 0
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_405
timestamp 0
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_417
timestamp 0
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_429
timestamp 0
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_441
timestamp 0
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_447
timestamp 0
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_449
timestamp 0
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_461
timestamp 0
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_473
timestamp 0
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_485
timestamp 0
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_497
timestamp 0
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_503
timestamp 0
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_505
timestamp 0
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_517
timestamp 0
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_529
timestamp 0
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_541
timestamp 0
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_553
timestamp 0
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_559
timestamp 0
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_561
timestamp 0
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_573
timestamp 0
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_585
timestamp 0
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_597
timestamp 0
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_609
timestamp 0
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_615
timestamp 0
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_89_617
timestamp 0
transform 1 0 57868 0 -1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_3
timestamp 0
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_15
timestamp 0
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_27
timestamp 0
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_29
timestamp 0
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_41
timestamp 0
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_53
timestamp 0
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_65
timestamp 0
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_77
timestamp 0
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_83
timestamp 0
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_85
timestamp 0
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_97
timestamp 0
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_109
timestamp 0
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_121
timestamp 0
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_133
timestamp 0
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_139
timestamp 0
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_141
timestamp 0
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_153
timestamp 0
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_165
timestamp 0
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_177
timestamp 0
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_189
timestamp 0
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_195
timestamp 0
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_197
timestamp 0
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_209
timestamp 0
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_221
timestamp 0
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_233
timestamp 0
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_245
timestamp 0
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_251
timestamp 0
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_253
timestamp 0
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_265
timestamp 0
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_277
timestamp 0
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_289
timestamp 0
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_301
timestamp 0
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_307
timestamp 0
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_309
timestamp 0
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_321
timestamp 0
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_333
timestamp 0
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_345
timestamp 0
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_357
timestamp 0
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_363
timestamp 0
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_365
timestamp 0
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_377
timestamp 0
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_389
timestamp 0
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_401
timestamp 0
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_413
timestamp 0
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_419
timestamp 0
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_421
timestamp 0
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_433
timestamp 0
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_445
timestamp 0
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_457
timestamp 0
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_469
timestamp 0
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_475
timestamp 0
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_477
timestamp 0
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_489
timestamp 0
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_501
timestamp 0
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_513
timestamp 0
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_525
timestamp 0
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_531
timestamp 0
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_533
timestamp 0
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_545
timestamp 0
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_557
timestamp 0
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_569
timestamp 0
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_581
timestamp 0
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_587
timestamp 0
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_589
timestamp 0
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_601
timestamp 0
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_613
timestamp 0
transform 1 0 57500 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_3
timestamp 0
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_15
timestamp 0
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_27
timestamp 0
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_39
timestamp 0
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91_51
timestamp 0
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_55
timestamp 0
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_57
timestamp 0
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_69
timestamp 0
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_81
timestamp 0
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_93
timestamp 0
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_105
timestamp 0
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_111
timestamp 0
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_113
timestamp 0
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_125
timestamp 0
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_137
timestamp 0
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_149
timestamp 0
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_161
timestamp 0
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_167
timestamp 0
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_169
timestamp 0
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_181
timestamp 0
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_193
timestamp 0
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_205
timestamp 0
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_217
timestamp 0
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_223
timestamp 0
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_225
timestamp 0
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_237
timestamp 0
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_249
timestamp 0
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_261
timestamp 0
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_273
timestamp 0
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_279
timestamp 0
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_281
timestamp 0
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_293
timestamp 0
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_305
timestamp 0
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_317
timestamp 0
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_329
timestamp 0
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_335
timestamp 0
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_337
timestamp 0
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_349
timestamp 0
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_361
timestamp 0
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_373
timestamp 0
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_385
timestamp 0
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_391
timestamp 0
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_393
timestamp 0
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_405
timestamp 0
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_417
timestamp 0
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_429
timestamp 0
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_441
timestamp 0
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_447
timestamp 0
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_449
timestamp 0
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_461
timestamp 0
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_473
timestamp 0
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_485
timestamp 0
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_497
timestamp 0
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_503
timestamp 0
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_505
timestamp 0
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_517
timestamp 0
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_529
timestamp 0
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_541
timestamp 0
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_553
timestamp 0
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_559
timestamp 0
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_561
timestamp 0
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_573
timestamp 0
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_585
timestamp 0
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_597
timestamp 0
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_609
timestamp 0
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_615
timestamp 0
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_91_617
timestamp 0
transform 1 0 57868 0 -1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_3
timestamp 0
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_15
timestamp 0
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_27
timestamp 0
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_29
timestamp 0
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_41
timestamp 0
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_53
timestamp 0
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_65
timestamp 0
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_77
timestamp 0
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_83
timestamp 0
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_85
timestamp 0
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_97
timestamp 0
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_109
timestamp 0
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_121
timestamp 0
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_133
timestamp 0
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_139
timestamp 0
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_141
timestamp 0
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_153
timestamp 0
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_165
timestamp 0
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_177
timestamp 0
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_189
timestamp 0
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_195
timestamp 0
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_197
timestamp 0
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_209
timestamp 0
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_221
timestamp 0
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_233
timestamp 0
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_245
timestamp 0
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_251
timestamp 0
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_253
timestamp 0
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_265
timestamp 0
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_277
timestamp 0
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_289
timestamp 0
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_301
timestamp 0
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_307
timestamp 0
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_309
timestamp 0
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_321
timestamp 0
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_333
timestamp 0
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_345
timestamp 0
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_357
timestamp 0
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_363
timestamp 0
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_365
timestamp 0
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_377
timestamp 0
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_389
timestamp 0
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_401
timestamp 0
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_413
timestamp 0
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_419
timestamp 0
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_421
timestamp 0
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_433
timestamp 0
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_445
timestamp 0
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_457
timestamp 0
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_469
timestamp 0
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_475
timestamp 0
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_477
timestamp 0
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_489
timestamp 0
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_501
timestamp 0
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_513
timestamp 0
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_525
timestamp 0
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_531
timestamp 0
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_533
timestamp 0
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_545
timestamp 0
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_557
timestamp 0
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_569
timestamp 0
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_581
timestamp 0
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_587
timestamp 0
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_589
timestamp 0
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_601
timestamp 0
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_613
timestamp 0
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_3
timestamp 0
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_15
timestamp 0
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_27
timestamp 0
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_39
timestamp 0
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93_51
timestamp 0
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_55
timestamp 0
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_57
timestamp 0
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_69
timestamp 0
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_81
timestamp 0
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_93
timestamp 0
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_105
timestamp 0
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_111
timestamp 0
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_113
timestamp 0
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_125
timestamp 0
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_137
timestamp 0
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_149
timestamp 0
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_161
timestamp 0
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_167
timestamp 0
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_169
timestamp 0
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_181
timestamp 0
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_93_193
timestamp 0
transform 1 0 18860 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_93_221
timestamp 0
transform 1 0 21436 0 -1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_225
timestamp 0
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_237
timestamp 0
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_249
timestamp 0
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_261
timestamp 0
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_273
timestamp 0
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_279
timestamp 0
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_281
timestamp 0
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_293
timestamp 0
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_305
timestamp 0
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_317
timestamp 0
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_329
timestamp 0
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_335
timestamp 0
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_337
timestamp 0
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_349
timestamp 0
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_361
timestamp 0
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_373
timestamp 0
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_385
timestamp 0
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_391
timestamp 0
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_393
timestamp 0
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_405
timestamp 0
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_417
timestamp 0
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_429
timestamp 0
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_441
timestamp 0
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_447
timestamp 0
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_449
timestamp 0
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_461
timestamp 0
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_473
timestamp 0
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_485
timestamp 0
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_497
timestamp 0
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_503
timestamp 0
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_505
timestamp 0
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_517
timestamp 0
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_529
timestamp 0
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_541
timestamp 0
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_553
timestamp 0
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_559
timestamp 0
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_561
timestamp 0
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_573
timestamp 0
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_585
timestamp 0
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_597
timestamp 0
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_609
timestamp 0
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_615
timestamp 0
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_93_617
timestamp 0
transform 1 0 57868 0 -1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_3
timestamp 0
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_15
timestamp 0
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_27
timestamp 0
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_29
timestamp 0
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_41
timestamp 0
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_53
timestamp 0
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_65
timestamp 0
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_77
timestamp 0
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_83
timestamp 0
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_85
timestamp 0
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_97
timestamp 0
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_109
timestamp 0
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_121
timestamp 0
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_133
timestamp 0
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_139
timestamp 0
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_141
timestamp 0
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_153
timestamp 0
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_165
timestamp 0
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_177
timestamp 0
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_189
timestamp 0
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_195
timestamp 0
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_197
timestamp 0
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94_209
timestamp 0
transform 1 0 20332 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_233
timestamp 0
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_245
timestamp 0
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_251
timestamp 0
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_253
timestamp 0
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_265
timestamp 0
transform 1 0 25484 0 1 53312
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_291
timestamp 0
transform 1 0 27876 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94_303
timestamp 0
transform 1 0 28980 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_307
timestamp 0
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_309
timestamp 0
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_321
timestamp 0
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_333
timestamp 0
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_345
timestamp 0
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_357
timestamp 0
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_363
timestamp 0
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_365
timestamp 0
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_377
timestamp 0
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_389
timestamp 0
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_401
timestamp 0
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_413
timestamp 0
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_419
timestamp 0
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_421
timestamp 0
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_433
timestamp 0
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_445
timestamp 0
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_457
timestamp 0
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_469
timestamp 0
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_475
timestamp 0
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_477
timestamp 0
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_489
timestamp 0
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_501
timestamp 0
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_513
timestamp 0
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_525
timestamp 0
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_531
timestamp 0
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_533
timestamp 0
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_545
timestamp 0
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_557
timestamp 0
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_569
timestamp 0
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_581
timestamp 0
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_587
timestamp 0
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_589
timestamp 0
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_601
timestamp 0
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_613
timestamp 0
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_3
timestamp 0
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_15
timestamp 0
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_27
timestamp 0
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_39
timestamp 0
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95_51
timestamp 0
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_55
timestamp 0
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_57
timestamp 0
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_69
timestamp 0
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_81
timestamp 0
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_93
timestamp 0
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_105
timestamp 0
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_111
timestamp 0
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_113
timestamp 0
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_125
timestamp 0
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_137
timestamp 0
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_149
timestamp 0
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_161
timestamp 0
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_167
timestamp 0
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_169
timestamp 0
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_181
timestamp 0
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_95_193
timestamp 0
transform 1 0 18860 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_95_201
timestamp 0
transform 1 0 19596 0 -1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_225
timestamp 0
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_237
timestamp 0
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_249
timestamp 0
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_261
timestamp 0
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_273
timestamp 0
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_279
timestamp 0
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_281
timestamp 0
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_293
timestamp 0
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_305
timestamp 0
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_317
timestamp 0
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_329
timestamp 0
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_335
timestamp 0
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_337
timestamp 0
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_349
timestamp 0
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_361
timestamp 0
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_373
timestamp 0
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_385
timestamp 0
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_391
timestamp 0
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_393
timestamp 0
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_405
timestamp 0
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_417
timestamp 0
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_429
timestamp 0
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_441
timestamp 0
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_447
timestamp 0
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_449
timestamp 0
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_461
timestamp 0
transform 1 0 43516 0 -1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_487
timestamp 0
transform 1 0 45908 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95_499
timestamp 0
transform 1 0 47012 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_503
timestamp 0
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_505
timestamp 0
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_517
timestamp 0
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_529
timestamp 0
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_541
timestamp 0
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_553
timestamp 0
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_559
timestamp 0
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_561
timestamp 0
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_573
timestamp 0
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_585
timestamp 0
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_597
timestamp 0
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_609
timestamp 0
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_615
timestamp 0
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_95_617
timestamp 0
transform 1 0 57868 0 -1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_3
timestamp 0
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_15
timestamp 0
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_27
timestamp 0
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_29
timestamp 0
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_41
timestamp 0
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_53
timestamp 0
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_65
timestamp 0
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_77
timestamp 0
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_83
timestamp 0
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_85
timestamp 0
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_97
timestamp 0
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_109
timestamp 0
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_121
timestamp 0
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_133
timestamp 0
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_139
timestamp 0
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_141
timestamp 0
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_153
timestamp 0
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_165
timestamp 0
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_177
timestamp 0
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_189
timestamp 0
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_195
timestamp 0
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_197
timestamp 0
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_96_209
timestamp 0
transform 1 0 20332 0 1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_253
timestamp 0
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_96_265
timestamp 0
transform 1 0 25484 0 1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_309
timestamp 0
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_321
timestamp 0
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_333
timestamp 0
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_345
timestamp 0
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_357
timestamp 0
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_363
timestamp 0
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_365
timestamp 0
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96_377
timestamp 0
transform 1 0 35788 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_381
timestamp 0
transform 1 0 36156 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_402
timestamp 0
transform 1 0 38088 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_414
timestamp 0
transform 1 0 39192 0 1 54400
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_461
timestamp 0
transform 1 0 43516 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_96_473
timestamp 0
transform 1 0 44620 0 1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_497
timestamp 0
transform 1 0 46828 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_509
timestamp 0
transform 1 0 47932 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_96_521
timestamp 0
transform 1 0 49036 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_96_529
timestamp 0
transform 1 0 49772 0 1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_533
timestamp 0
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_545
timestamp 0
transform 1 0 51244 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_572
timestamp 0
transform 1 0 53728 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_96_584
timestamp 0
transform 1 0 54832 0 1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_589
timestamp 0
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_601
timestamp 0
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_613
timestamp 0
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_3
timestamp 0
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_15
timestamp 0
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_27
timestamp 0
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_39
timestamp 0
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97_51
timestamp 0
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_55
timestamp 0
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_57
timestamp 0
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_69
timestamp 0
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_81
timestamp 0
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_93
timestamp 0
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_105
timestamp 0
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_111
timestamp 0
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_113
timestamp 0
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_125
timestamp 0
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_137
timestamp 0
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_149
timestamp 0
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_161
timestamp 0
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_167
timestamp 0
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_97_175
timestamp 0
transform 1 0 17204 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_97_181
timestamp 0
transform 1 0 17756 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97_233
timestamp 0
transform 1 0 22540 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_97_277
timestamp 0
transform 1 0 26588 0 -1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_281
timestamp 0
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_293
timestamp 0
transform 1 0 28060 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_314
timestamp 0
transform 1 0 29992 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97_326
timestamp 0
transform 1 0 31096 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_97_334
timestamp 0
transform 1 0 31832 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_377
timestamp 0
transform 1 0 35788 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_97_389
timestamp 0
transform 1 0 36892 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97_393
timestamp 0
transform 1 0 37260 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_441
timestamp 0
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_447
timestamp 0
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_449
timestamp 0
transform 1 0 42412 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97_495
timestamp 0
transform 1 0 46644 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_503
timestamp 0
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_505
timestamp 0
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_97_517
timestamp 0
transform 1 0 48668 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_539
timestamp 0
transform 1 0 50692 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_581
timestamp 0
transform 1 0 54556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_593
timestamp 0
transform 1 0 55660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97_605
timestamp 0
transform 1 0 56764 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_97_613
timestamp 0
transform 1 0 57500 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97_617
timestamp 0
transform 1 0 57868 0 -1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_3
timestamp 0
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_15
timestamp 0
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_27
timestamp 0
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_29
timestamp 0
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_41
timestamp 0
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_53
timestamp 0
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_65
timestamp 0
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_77
timestamp 0
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_83
timestamp 0
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_85
timestamp 0
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_97
timestamp 0
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_109
timestamp 0
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_121
timestamp 0
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_133
timestamp 0
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_139
timestamp 0
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_141
timestamp 0
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_153
timestamp 0
transform 1 0 15180 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_186
timestamp 0
transform 1 0 18216 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_98_190
timestamp 0
transform 1 0 18584 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_205
timestamp 0
transform 1 0 19964 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_211
timestamp 0
transform 1 0 20516 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_259
timestamp 0
transform 1 0 24932 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_98_271
timestamp 0
transform 1 0 26036 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_296
timestamp 0
transform 1 0 28336 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_317
timestamp 0
transform 1 0 30268 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_329
timestamp 0
transform 1 0 31372 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_341
timestamp 0
transform 1 0 32476 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_98_353
timestamp 0
transform 1 0 33580 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_98_361
timestamp 0
transform 1 0 34316 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_98_365
timestamp 0
transform 1 0 34684 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_369
timestamp 0
transform 1 0 35052 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_376
timestamp 0
transform 1 0 35696 0 1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_402
timestamp 0
transform 1 0 38088 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_414
timestamp 0
transform 1 0 39192 0 1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_421
timestamp 0
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_433
timestamp 0
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_445
timestamp 0
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_457
timestamp 0
transform 1 0 43148 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_461
timestamp 0
transform 1 0 43516 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_485
timestamp 0
transform 1 0 45724 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_497
timestamp 0
transform 1 0 46828 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_509
timestamp 0
transform 1 0 47932 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_98_521
timestamp 0
transform 1 0 49036 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_98_529
timestamp 0
transform 1 0 49772 0 1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_533
timestamp 0
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_545
timestamp 0
transform 1 0 51244 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_566
timestamp 0
transform 1 0 53176 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_98_578
timestamp 0
transform 1 0 54280 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_98_586
timestamp 0
transform 1 0 55016 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_589
timestamp 0
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_601
timestamp 0
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_613
timestamp 0
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_3
timestamp 0
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_15
timestamp 0
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_27
timestamp 0
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_39
timestamp 0
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99_51
timestamp 0
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_55
timestamp 0
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_57
timestamp 0
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_69
timestamp 0
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_81
timestamp 0
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_93
timestamp 0
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_105
timestamp 0
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_111
timestamp 0
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_113
timestamp 0
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_125
timestamp 0
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_137
timestamp 0
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_149
timestamp 0
transform 1 0 14812 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99_169
timestamp 0
transform 1 0 16652 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_99_237
timestamp 0
transform 1 0 22908 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_252
timestamp 0
transform 1 0 24288 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_270
timestamp 0
transform 1 0 25944 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99_284
timestamp 0
transform 1 0 27232 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_304
timestamp 0
transform 1 0 29072 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_316
timestamp 0
transform 1 0 30176 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99_328
timestamp 0
transform 1 0 31280 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_332
timestamp 0
transform 1 0 31648 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_99_346
timestamp 0
transform 1 0 32936 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_99_354
timestamp 0
transform 1 0 33672 0 -1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_369
timestamp 0
transform 1 0 35052 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99_381
timestamp 0
transform 1 0 36156 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_396
timestamp 0
transform 1 0 37536 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99_414
timestamp 0
transform 1 0 39192 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_99_430
timestamp 0
transform 1 0 40664 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_438
timestamp 0
transform 1 0 41400 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_442
timestamp 0
transform 1 0 41768 0 -1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_485
timestamp 0
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_497
timestamp 0
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_503
timestamp 0
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_505
timestamp 0
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_99_517
timestamp 0
transform 1 0 48668 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_99_532
timestamp 0
transform 1 0 50048 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99_558
timestamp 0
transform 1 0 52440 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_578
timestamp 0
transform 1 0 54280 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_590
timestamp 0
transform 1 0 55384 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_602
timestamp 0
transform 1 0 56488 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99_614
timestamp 0
transform 1 0 57592 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_99_617
timestamp 0
transform 1 0 57868 0 -1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_3
timestamp 0
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_15
timestamp 0
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_27
timestamp 0
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_29
timestamp 0
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_41
timestamp 0
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_53
timestamp 0
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_65
timestamp 0
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_77
timestamp 0
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_83
timestamp 0
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_85
timestamp 0
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_97
timestamp 0
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_109
timestamp 0
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_121
timestamp 0
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_133
timestamp 0
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_139
timestamp 0
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_141
timestamp 0
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100_153
timestamp 0
transform 1 0 15180 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_190
timestamp 0
transform 1 0 18584 0 1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_197
timestamp 0
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_209
timestamp 0
transform 1 0 20332 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_100_230
timestamp 0
transform 1 0 22264 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_246
timestamp 0
transform 1 0 23736 0 1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_253
timestamp 0
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_100_265
timestamp 0
transform 1 0 25484 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100_273
timestamp 0
transform 1 0 26220 0 1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_295
timestamp 0
transform 1 0 28244 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_307
timestamp 0
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_309
timestamp 0
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_321
timestamp 0
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_333
timestamp 0
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_345
timestamp 0
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_357
timestamp 0
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_363
timestamp 0
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_365
timestamp 0
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_377
timestamp 0
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_389
timestamp 0
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_401
timestamp 0
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_413
timestamp 0
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_419
timestamp 0
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_421
timestamp 0
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_433
timestamp 0
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_445
timestamp 0
transform 1 0 42044 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_457
timestamp 0
transform 1 0 43148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_469
timestamp 0
transform 1 0 44252 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_475
timestamp 0
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_477
timestamp 0
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_489
timestamp 0
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_501
timestamp 0
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_513
timestamp 0
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_525
timestamp 0
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_531
timestamp 0
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_533
timestamp 0
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100_545
timestamp 0
transform 1 0 51244 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_568
timestamp 0
transform 1 0 53360 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_100_580
timestamp 0
transform 1 0 54464 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_589
timestamp 0
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_601
timestamp 0
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_613
timestamp 0
transform 1 0 57500 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_101_13
timestamp 0
transform 1 0 2300 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_19
timestamp 0
transform 1 0 2852 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_101_26
timestamp 0
transform 1 0 3496 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_29
timestamp 0
transform 1 0 3772 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101_47
timestamp 0
transform 1 0 5428 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_55
timestamp 0
transform 1 0 6164 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_57
timestamp 0
transform 1 0 6348 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_61
timestamp 0
transform 1 0 6716 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_68
timestamp 0
transform 1 0 7360 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_80
timestamp 0
transform 1 0 8464 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_91
timestamp 0
transform 1 0 9476 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_103
timestamp 0
transform 1 0 10580 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_101_110
timestamp 0
transform 1 0 11224 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_113
timestamp 0
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101_131
timestamp 0
transform 1 0 13156 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_139
timestamp 0
transform 1 0 13892 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_141
timestamp 0
transform 1 0 14076 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_145
timestamp 0
transform 1 0 14444 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_152
timestamp 0
transform 1 0 15088 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_164
timestamp 0
transform 1 0 16192 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_175
timestamp 0
transform 1 0 17204 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_187
timestamp 0
transform 1 0 18308 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_101_194
timestamp 0
transform 1 0 18952 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_197
timestamp 0
transform 1 0 19228 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101_215
timestamp 0
transform 1 0 20884 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_223
timestamp 0
transform 1 0 21620 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_225
timestamp 0
transform 1 0 21804 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_229
timestamp 0
transform 1 0 22172 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_236
timestamp 0
transform 1 0 22816 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_248
timestamp 0
transform 1 0 23920 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_259
timestamp 0
transform 1 0 24932 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_271
timestamp 0
transform 1 0 26036 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_101_278
timestamp 0
transform 1 0 26680 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_281
timestamp 0
transform 1 0 26956 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101_299
timestamp 0
transform 1 0 28612 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_307
timestamp 0
transform 1 0 29348 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_309
timestamp 0
transform 1 0 29532 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_313
timestamp 0
transform 1 0 29900 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_320
timestamp 0
transform 1 0 30544 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_332
timestamp 0
transform 1 0 31648 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_343
timestamp 0
transform 1 0 32660 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_355
timestamp 0
transform 1 0 33764 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_101_362
timestamp 0
transform 1 0 34408 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_365
timestamp 0
transform 1 0 34684 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101_383
timestamp 0
transform 1 0 36340 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_391
timestamp 0
transform 1 0 37076 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_393
timestamp 0
transform 1 0 37260 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_397
timestamp 0
transform 1 0 37628 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_404
timestamp 0
transform 1 0 38272 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_416
timestamp 0
transform 1 0 39376 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_427
timestamp 0
transform 1 0 40388 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_439
timestamp 0
transform 1 0 41492 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_101_446
timestamp 0
transform 1 0 42136 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_449
timestamp 0
transform 1 0 42412 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101_467
timestamp 0
transform 1 0 44068 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_475
timestamp 0
transform 1 0 44804 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_477
timestamp 0
transform 1 0 44988 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_481
timestamp 0
transform 1 0 45356 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_488
timestamp 0
transform 1 0 46000 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_500
timestamp 0
transform 1 0 47104 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_511
timestamp 0
transform 1 0 48116 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_523
timestamp 0
transform 1 0 49220 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_101_530
timestamp 0
transform 1 0 49864 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_533
timestamp 0
transform 1 0 50140 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101_551
timestamp 0
transform 1 0 51796 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_559
timestamp 0
transform 1 0 52532 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_561
timestamp 0
transform 1 0 52716 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_565
timestamp 0
transform 1 0 53084 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_572
timestamp 0
transform 1 0 53728 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_584
timestamp 0
transform 1 0 54832 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_595
timestamp 0
transform 1 0 55844 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_607
timestamp 0
transform 1 0 56948 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_101_614
timestamp 0
transform 1 0 57592 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_101_617
timestamp 0
transform 1 0 57868 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 0
transform -1 0 30268 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 0
transform -1 0 45724 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 0
transform 1 0 21804 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 0
transform -1 0 54280 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 0
transform -1 0 27232 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 0
transform -1 0 27968 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 0
transform -1 0 44344 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 0
transform 1 0 23000 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  input1
timestamp 0
transform -1 0 58604 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 0
transform 1 0 1380 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  output3
timestamp 0
transform -1 0 3496 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output4
timestamp 0
transform -1 0 22816 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output5
timestamp 0
transform -1 0 24932 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output6
timestamp 0
transform -1 0 26680 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output7
timestamp 0
transform 1 0 28060 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output8
timestamp 0
transform 1 0 29992 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output9
timestamp 0
transform -1 0 32660 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output10
timestamp 0
transform -1 0 34408 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output11
timestamp 0
transform -1 0 36340 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output12
timestamp 0
transform -1 0 38272 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output13
timestamp 0
transform -1 0 40388 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output14
timestamp 0
transform -1 0 5428 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output15
timestamp 0
transform -1 0 42136 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 0
transform -1 0 44068 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 0
transform 1 0 45448 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output18
timestamp 0
transform 1 0 47564 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output19
timestamp 0
transform 1 0 49312 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output20
timestamp 0
transform 1 0 51244 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 0
transform 1 0 53176 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 0
transform 1 0 55292 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 0
transform 1 0 57040 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 0
transform 1 0 58052 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 0
transform -1 0 7360 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 0
transform -1 0 9476 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 0
transform -1 0 11224 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output28
timestamp 0
transform -1 0 13156 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output29
timestamp 0
transform -1 0 15088 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 0
transform -1 0 17204 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output31
timestamp 0
transform -1 0 18952 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 0
transform -1 0 20884 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 0
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 0
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 0
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 0
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 0
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 0
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 0
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 0
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 0
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 0
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 0
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 0
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 0
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 0
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 0
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 0
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 0
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 0
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 0
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 0
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 0
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 0
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 0
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 0
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 0
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 0
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 0
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 0
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 0
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 0
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 0
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 0
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 0
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 0
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 0
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 0
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 0
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 0
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 0
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 0
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 0
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 0
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 0
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 0
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 0
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 0
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 0
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 0
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 0
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 0
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 0
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 0
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 0
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 0
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 0
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 0
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 0
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 0
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 0
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 0
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 0
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 0
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 0
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 0
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 0
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 0
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 0
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 0
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 0
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 0
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 0
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 0
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 0
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 0
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 0
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 0
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 0
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 0
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 0
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 0
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 0
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 0
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 0
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 0
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 0
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 0
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 0
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 0
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 0
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 0
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 0
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 0
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 0
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 0
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 0
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 0
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 0
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 0
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 0
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 0
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 0
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 0
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 0
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 0
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 0
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 0
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 0
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 0
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 0
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 0
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 0
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 0
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 0
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 0
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 0
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 0
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 0
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 0
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 0
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 0
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 0
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 0
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 0
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 0
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 0
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 0
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 0
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 0
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 0
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 0
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 0
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 0
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 0
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 0
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 0
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 0
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 0
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 0
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 0
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 0
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 0
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 0
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 0
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 0
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 0
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 0
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 0
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 0
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 0
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 0
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 0
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 0
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 0
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 0
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 0
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 0
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 0
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 0
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 0
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 0
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 0
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 0
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 0
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 0
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 0
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 0
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 0
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 0
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 0
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 0
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 0
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 0
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 0
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 0
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 0
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 0
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 0
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 0
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 0
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 0
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 0
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 0
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 0
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 0
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 0
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 0
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 0
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 0
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 0
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 0
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 0
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 0
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 0
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 0
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 0
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 0
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 0
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 0
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 0
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 0
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 0
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 0
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 0
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 0
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 0
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 0
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 0
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 0
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 0
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 0
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 0
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 0
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 0
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 0
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 0
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 0
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 0
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 0
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 0
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 0
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 0
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 0
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 0
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 0
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 0
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 0
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 0
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 0
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 0
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 0
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 0
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 0
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 0
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 0
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 0
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 0
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 0
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 0
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 0
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 0
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 0
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 0
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 0
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 0
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 0
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 0
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 0
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 0
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 0
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 0
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 0
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 0
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 0
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 0
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 0
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 0
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 0
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 0
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 0
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 0
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 0
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 0
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 0
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 0
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 0
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 0
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 0
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 0
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 0
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 0
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 0
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 0
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 0
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 0
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 0
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 0
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 0
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 0
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 0
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 0
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 0
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 0
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 0
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 0
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 0
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 0
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 0
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 0
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 0
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 0
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 0
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 0
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 0
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 0
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 0
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 0
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 0
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 0
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 0
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 0
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 0
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 0
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 0
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 0
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 0
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 0
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 0
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 0
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 0
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 0
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 0
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 0
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 0
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 0
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 0
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 0
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 0
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 0
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 0
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 0
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 0
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 0
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 0
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 0
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 0
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 0
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 0
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 0
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 0
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 0
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 0
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 0
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 0
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 0
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 0
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 0
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 0
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 0
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 0
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 0
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 0
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 0
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 0
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 0
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 0
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 0
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 0
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 0
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 0
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 0
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 0
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 0
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 0
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 0
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 0
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 0
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 0
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 0
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 0
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 0
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 0
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 0
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 0
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 0
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 0
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 0
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 0
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 0
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 0
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 0
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 0
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 0
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 0
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 0
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 0
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 0
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 0
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 0
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 0
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 0
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 0
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 0
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 0
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 0
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 0
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 0
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 0
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 0
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 0
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 0
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 0
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 0
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 0
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 0
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 0
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 0
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 0
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 0
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 0
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 0
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 0
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 0
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 0
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 0
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 0
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 0
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 0
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 0
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 0
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 0
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 0
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 0
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 0
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 0
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 0
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 0
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 0
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 0
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 0
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 0
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 0
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 0
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 0
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 0
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 0
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 0
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 0
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 0
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 0
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 0
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 0
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 0
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 0
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 0
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 0
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 0
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 0
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 0
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 0
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 0
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 0
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 0
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 0
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 0
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 0
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 0
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 0
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 0
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 0
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 0
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 0
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 0
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 0
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 0
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 0
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 0
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 0
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 0
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 0
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 0
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 0
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 0
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 0
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 0
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 0
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 0
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 0
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 0
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 0
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 0
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 0
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 0
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 0
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 0
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 0
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 0
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 0
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 0
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 0
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 0
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 0
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 0
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 0
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 0
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 0
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 0
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 0
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 0
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 0
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 0
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 0
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 0
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 0
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 0
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 0
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 0
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 0
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 0
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 0
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 0
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 0
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 0
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 0
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 0
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 0
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 0
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 0
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 0
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 0
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 0
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 0
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 0
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 0
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 0
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 0
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 0
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 0
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 0
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 0
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 0
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 0
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 0
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 0
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 0
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 0
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 0
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 0
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 0
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 0
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 0
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 0
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 0
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 0
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 0
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 0
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 0
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 0
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 0
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 0
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 0
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 0
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 0
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 0
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 0
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 0
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 0
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 0
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 0
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 0
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 0
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 0
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 0
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 0
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 0
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 0
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 0
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 0
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 0
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 0
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 0
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 0
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 0
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 0
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 0
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 0
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 0
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 0
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 0
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 0
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 0
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 0
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 0
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 0
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 0
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 0
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 0
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 0
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 0
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 0
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 0
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 0
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 0
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 0
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 0
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 0
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 0
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 0
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 0
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 0
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 0
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 0
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 0
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 0
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 0
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 0
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 0
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 0
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 0
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 0
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 0
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 0
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 0
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 0
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 0
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 0
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 0
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 0
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 0
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 0
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 0
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 0
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 0
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 0
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 0
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 0
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 0
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 0
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 0
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 0
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 0
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 0
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 0
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 0
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 0
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 0
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 0
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 0
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 0
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 0
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 0
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 0
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 0
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 0
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 0
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 0
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 0
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 0
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 0
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 0
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 0
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 0
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 0
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 0
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 0
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 0
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 0
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 0
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 0
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 0
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 0
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 0
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 0
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 0
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 0
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 0
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 0
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 0
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 0
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 0
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 0
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 0
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 0
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 0
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 0
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 0
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 0
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 0
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 0
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 0
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 0
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 0
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 0
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 0
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 0
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 0
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 0
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 0
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 0
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 0
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 0
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 0
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 0
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 0
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 0
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 0
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 0
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 0
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 0
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 0
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 0
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 0
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 0
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 0
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 0
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 0
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 0
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 0
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 0
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 0
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 0
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 0
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 0
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 0
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 0
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 0
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 0
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 0
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 0
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 0
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 0
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 0
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 0
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 0
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 0
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 0
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 0
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 0
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 0
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 0
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 0
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 0
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 0
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 0
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 0
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 0
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 0
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 0
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 0
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 0
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 0
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 0
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 0
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 0
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 0
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 0
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 0
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 0
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 0
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 0
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 0
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 0
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 0
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 0
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 0
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 0
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 0
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 0
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 0
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 0
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 0
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 0
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 0
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 0
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 0
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 0
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 0
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 0
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 0
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 0
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 0
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 0
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 0
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 0
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 0
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 0
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 0
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 0
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 0
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 0
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 0
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 0
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 0
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 0
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 0
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 0
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 0
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 0
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 0
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 0
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 0
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 0
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 0
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 0
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 0
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 0
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 0
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 0
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 0
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 0
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 0
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 0
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 0
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 0
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 0
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 0
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 0
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 0
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 0
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 0
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 0
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 0
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 0
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 0
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 0
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 0
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 0
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 0
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 0
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 0
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 0
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 0
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 0
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 0
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 0
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 0
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 0
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 0
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 0
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 0
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 0
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 0
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 0
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 0
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 0
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 0
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 0
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 0
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 0
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 0
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 0
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 0
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 0
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 0
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 0
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 0
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 0
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 0
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 0
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 0
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 0
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 0
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 0
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 0
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 0
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 0
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 0
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 0
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 0
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 0
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 0
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 0
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 0
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 0
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 0
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 0
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 0
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 0
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 0
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 0
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 0
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 0
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 0
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 0
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 0
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 0
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 0
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 0
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 0
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 0
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 0
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 0
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 0
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 0
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 0
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 0
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 0
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 0
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 0
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 0
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 0
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 0
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 0
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 0
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 0
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 0
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 0
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 0
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 0
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 0
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 0
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 0
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 0
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 0
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 0
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 0
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 0
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 0
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 0
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 0
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 0
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 0
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 0
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 0
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 0
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 0
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 0
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 0
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 0
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 0
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 0
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 0
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 0
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 0
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 0
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 0
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 0
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 0
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 0
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 0
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 0
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 0
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 0
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 0
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 0
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 0
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 0
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 0
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 0
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 0
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 0
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 0
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 0
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 0
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 0
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 0
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 0
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 0
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 0
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 0
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 0
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 0
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 0
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 0
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 0
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 0
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 0
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 0
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 0
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 0
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 0
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 0
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 0
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 0
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 0
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 0
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 0
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 0
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 0
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 0
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 0
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 0
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 0
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 0
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 0
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 0
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 0
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 0
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 0
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 0
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 0
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 0
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 0
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 0
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 0
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 0
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 0
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 0
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 0
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 0
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 0
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 0
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 0
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 0
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 0
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 0
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 0
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 0
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 0
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 0
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 0
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 0
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 0
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 0
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 0
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 0
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 0
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 0
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 0
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 0
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 0
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 0
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 0
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 0
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 0
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 0
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 0
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 0
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 0
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 0
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 0
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 0
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 0
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 0
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 0
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 0
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 0
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 0
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 0
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 0
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 0
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 0
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 0
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 0
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 0
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 0
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 0
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 0
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 0
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 0
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 0
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 0
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 0
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 0
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 0
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 0
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 0
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 0
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 0
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 0
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 0
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 0
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 0
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 0
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 0
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 0
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 0
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 0
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 0
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 0
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 0
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 0
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 0
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 0
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 0
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 0
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 0
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 0
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 0
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 0
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 0
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 0
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 0
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 0
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 0
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 0
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 0
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 0
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 0
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 0
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 0
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 0
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 0
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 0
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 0
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 0
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 0
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 0
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 0
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 0
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 0
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 0
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 0
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 0
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 0
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 0
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 0
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 0
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 0
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 0
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 0
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 0
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 0
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 0
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 0
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 0
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 0
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 0
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 0
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 0
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 0
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 0
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 0
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 0
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 0
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 0
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 0
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 0
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 0
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 0
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 0
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 0
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 0
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 0
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 0
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 0
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 0
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 0
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 0
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 0
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 0
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 0
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 0
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 0
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 0
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 0
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 0
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 0
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 0
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 0
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 0
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 0
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 0
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 0
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 0
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 0
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 0
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 0
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 0
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 0
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 0
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 0
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 0
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 0
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 0
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 0
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 0
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 0
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 0
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 0
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 0
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 0
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 0
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 0
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 0
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 0
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 0
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 0
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 0
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 0
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 0
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 0
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 0
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 0
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 0
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 0
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 0
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 0
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 0
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 0
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 0
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 0
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 0
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 0
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 0
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 0
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 0
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 0
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 0
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 0
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 0
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 0
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 0
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 0
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 0
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 0
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 0
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 0
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 0
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 0
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 0
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 0
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 0
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 0
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 0
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 0
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 0
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 0
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 0
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 0
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 0
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 0
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 0
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 0
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 0
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 0
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 0
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 0
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 0
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 0
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 0
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 0
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 0
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 0
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 0
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 0
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 0
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 0
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 0
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 0
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 0
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 0
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 0
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 0
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 0
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 0
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 0
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 0
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 0
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 0
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 0
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 0
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 0
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 0
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 0
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 0
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 0
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 0
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 0
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 0
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 0
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 0
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 0
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 0
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 0
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 0
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 0
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 0
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 0
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 0
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 0
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 0
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 0
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 0
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 0
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 0
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
<< labels >>
rlabel metal1 s 29992 57664 29992 57664 4 VGND
rlabel metal1 s 29992 57120 29992 57120 4 VPWR
rlabel metal2 s 32430 55726 32430 55726 4 _000_
rlabel metal1 s 34546 55182 34546 55182 4 _001_
rlabel metal1 s 37628 56134 37628 56134 4 _002_
rlabel metal2 s 38663 55284 38663 55284 4 _003_
rlabel metal1 s 39974 56134 39974 56134 4 _004_
rlabel metal1 s 41860 56134 41860 56134 4 _005_
rlabel metal2 s 43286 55454 43286 55454 4 _006_
rlabel metal1 s 44850 55182 44850 55182 4 _007_
rlabel metal1 s 44528 54230 44528 54230 4 _008_
rlabel metal1 s 49496 55182 49496 55182 4 _009_
rlabel metal2 s 51106 55726 51106 55726 4 _010_
rlabel metal1 s 52118 56134 52118 56134 4 _011_
rlabel metal1 s 51382 56202 51382 56202 4 _012_
rlabel metal2 s 51658 56236 51658 56236 4 _013_
rlabel metal1 s 21298 55624 21298 55624 4 _014_
rlabel metal1 s 21344 56406 21344 56406 4 _015_
rlabel metal2 s 16790 55420 16790 55420 4 _016_
rlabel metal1 s 16790 56984 16790 56984 4 _017_
rlabel metal2 s 15962 55046 15962 55046 4 _018_
rlabel metal2 s 17894 56372 17894 56372 4 _019_
rlabel metal1 s 20654 56712 20654 56712 4 _020_
rlabel metal1 s 18722 55386 18722 55386 4 _021_
rlabel metal1 s 18952 55862 18952 55862 4 _022_
rlabel metal1 s 20286 55590 20286 55590 4 _023_
rlabel metal2 s 22402 56032 22402 56032 4 _024_
rlabel metal2 s 22770 55896 22770 55896 4 _025_
rlabel metal2 s 25070 55726 25070 55726 4 _026_
rlabel metal1 s 26772 55794 26772 55794 4 _027_
rlabel metal2 s 27922 55692 27922 55692 4 _028_
rlabel metal2 s 28474 55454 28474 55454 4 _029_
rlabel metal1 s 15732 55726 15732 55726 4 _030_
rlabel metal2 s 16054 55930 16054 55930 4 _031_
rlabel metal1 s 22034 56338 22034 56338 4 _032_
rlabel metal2 s 18170 56372 18170 56372 4 _033_
rlabel metal2 s 17526 55692 17526 55692 4 _034_
rlabel metal2 s 18354 55930 18354 55930 4 _035_
rlabel metal2 s 19734 55930 19734 55930 4 _036_
rlabel metal1 s 22724 56338 22724 56338 4 _037_
rlabel metal1 s 24104 56338 24104 56338 4 _038_
rlabel metal1 s 25898 56262 25898 56262 4 _039_
rlabel metal1 s 27324 56474 27324 56474 4 _040_
rlabel metal2 s 28198 56644 28198 56644 4 _041_
rlabel metal2 s 28106 55930 28106 55930 4 _042_
rlabel metal1 s 19458 55760 19458 55760 4 _043_
rlabel metal1 s 31970 56338 31970 56338 4 _044_
rlabel metal1 s 34960 56338 34960 56338 4 _045_
rlabel metal1 s 37260 56338 37260 56338 4 _046_
rlabel metal1 s 39008 56338 39008 56338 4 _047_
rlabel metal1 s 39744 56338 39744 56338 4 _048_
rlabel metal1 s 41998 56338 41998 56338 4 _049_
rlabel metal2 s 43470 55930 43470 55930 4 _050_
rlabel metal2 s 44390 55930 44390 55930 4 _051_
rlabel metal1 s 44896 55726 44896 55726 4 _052_
rlabel metal1 s 17250 55794 17250 55794 4 _053_
rlabel metal1 s 50002 56270 50002 56270 4 _054_
rlabel metal1 s 51980 56338 51980 56338 4 _055_
rlabel metal1 s 52440 56338 52440 56338 4 _056_
rlabel metal1 s 50968 56338 50968 56338 4 _057_
rlabel metal2 s 52762 56644 52762 56644 4 _058_
rlabel metal1 s 19090 55726 19090 55726 4 _059_
rlabel metal1 s 16652 55930 16652 55930 4 _060_
rlabel metal2 s 16974 56202 16974 56202 4 _061_
rlabel metal1 s 15732 56814 15732 56814 4 _062_
rlabel metal2 s 38042 30335 38042 30335 4 clk
rlabel metal1 s 36248 55658 36248 55658 4 clknet_0_clk
rlabel metal1 s 26266 54740 26266 54740 4 clknet_2_0__leaf_clk
rlabel metal1 s 21666 56236 21666 56236 4 clknet_2_1__leaf_clk
rlabel metal1 s 37996 55250 37996 55250 4 clknet_2_2__leaf_clk
rlabel metal1 s 44850 55318 44850 55318 4 clknet_2_3__leaf_clk
rlabel metal2 s 58282 49776 58282 49776 4 net1
rlabel metal2 s 34270 56848 34270 56848 4 net10
rlabel metal2 s 35926 55930 35926 55930 4 net11
rlabel metal1 s 36524 56338 36524 56338 4 net12
rlabel metal1 s 40296 56474 40296 56474 4 net13
rlabel metal2 s 5290 57188 5290 57188 4 net14
rlabel metal2 s 41630 55828 41630 55828 4 net15
rlabel metal1 s 44068 55726 44068 55726 4 net16
rlabel metal2 s 44758 55522 44758 55522 4 net17
rlabel metal1 s 44942 56406 44942 56406 4 net18
rlabel metal1 s 49358 56474 49358 56474 4 net19
rlabel metal1 s 16928 56406 16928 56406 4 net2
rlabel metal1 s 51290 56406 51290 56406 4 net20
rlabel metal2 s 52026 57154 52026 57154 4 net21
rlabel metal2 s 53038 57188 53038 57188 4 net22
rlabel metal2 s 55890 56916 55890 56916 4 net23
rlabel metal2 s 56166 56916 56166 56916 4 net24
rlabel metal1 s 17664 56746 17664 56746 4 net25
rlabel metal2 s 15226 56984 15226 56984 4 net26
rlabel metal1 s 16698 56406 16698 56406 4 net27
rlabel metal1 s 18170 55794 18170 55794 4 net28
rlabel metal1 s 17342 56474 17342 56474 4 net29
rlabel metal2 s 4094 56610 4094 56610 4 net3
rlabel metal2 s 18722 56100 18722 56100 4 net30
rlabel metal1 s 19688 56270 19688 56270 4 net31
rlabel metal1 s 19734 56202 19734 56202 4 net32
rlabel metal1 s 29164 55862 29164 55862 4 net33
rlabel metal1 s 44712 56270 44712 56270 4 net34
rlabel metal1 s 22402 55250 22402 55250 4 net35
rlabel metal1 s 53360 56338 53360 56338 4 net36
rlabel metal1 s 26450 56474 26450 56474 4 net37
rlabel metal2 s 27186 56508 27186 56508 4 net38
rlabel metal1 s 43700 55930 43700 55930 4 net39
rlabel metal1 s 22356 56338 22356 56338 4 net4
rlabel metal1 s 23598 56474 23598 56474 4 net40
rlabel metal1 s 19373 55318 19373 55318 4 net41
rlabel metal1 s 35519 55318 35519 55318 4 net42
rlabel metal1 s 38035 55318 38035 55318 4 net43
rlabel metal1 s 24978 56474 24978 56474 4 net5
rlabel metal2 s 27094 56100 27094 56100 4 net6
rlabel metal2 s 27738 56916 27738 56916 4 net7
rlabel metal2 s 30130 56610 30130 56610 4 net8
rlabel metal1 s 32568 56474 32568 56474 4 net9
rlabel metal2 s 58558 44897 58558 44897 4 reset
rlabel metal1 s 1196 57426 1196 57426 4 scan_in
rlabel metal1 s 2944 57494 2944 57494 4 scan_out[0]
rlabel metal1 s 22264 57494 22264 57494 4 scan_out[10]
rlabel metal1 s 24288 57494 24288 57494 4 scan_out[11]
rlabel metal2 s 26266 57715 26266 57715 4 scan_out[12]
rlabel metal1 s 28152 57562 28152 57562 4 scan_out[13]
rlabel metal2 s 30406 57715 30406 57715 4 scan_out[14]
rlabel metal1 s 32016 57494 32016 57494 4 scan_out[15]
rlabel metal2 s 34178 58395 34178 58395 4 scan_out[16]
rlabel metal2 s 35742 58388 35742 58388 4 scan_out[17]
rlabel metal1 s 37720 57494 37720 57494 4 scan_out[18]
rlabel metal1 s 39744 57494 39744 57494 4 scan_out[19]
rlabel metal1 s 4876 57494 4876 57494 4 scan_out[1]
rlabel metal1 s 41584 57494 41584 57494 4 scan_out[20]
rlabel metal1 s 43516 57494 43516 57494 4 scan_out[21]
rlabel metal2 s 45402 58388 45402 58388 4 scan_out[22]
rlabel metal1 s 47564 57562 47564 57562 4 scan_out[23]
rlabel metal2 s 49680 57562 49680 57562 4 scan_out[24]
rlabel metal1 s 51336 57562 51336 57562 4 scan_out[25]
rlabel metal1 s 53268 57562 53268 57562 4 scan_out[26]
rlabel metal2 s 55062 58388 55062 58388 4 scan_out[27]
rlabel metal1 s 57132 57562 57132 57562 4 scan_out[28]
rlabel metal1 s 58742 57494 58742 57494 4 scan_out[29]
rlabel metal2 s 6762 58388 6762 58388 4 scan_out[2]
rlabel metal1 s 8832 57494 8832 57494 4 scan_out[3]
rlabel metal1 s 10672 57494 10672 57494 4 scan_out[4]
rlabel metal1 s 12604 57494 12604 57494 4 scan_out[5]
rlabel metal1 s 14536 57494 14536 57494 4 scan_out[6]
rlabel metal2 s 16422 58354 16422 58354 4 scan_out[7]
rlabel metal1 s 18400 57494 18400 57494 4 scan_out[8]
rlabel metal1 s 20332 57494 20332 57494 4 scan_out[9]
flabel metal5 s 1056 34712 58928 35032 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 4076 58928 4396 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 33724 2128 34044 57712 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 3004 2128 3324 57712 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 34052 58928 34372 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 3416 58928 3736 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 33064 2128 33384 57712 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 2344 2128 2664 57712 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 59200 14968 60000 15088 0 FreeSans 600 0 0 0 clk
port 3 nsew
flabel metal3 s 59200 44888 60000 45008 0 FreeSans 600 0 0 0 reset
port 4 nsew
flabel metal2 s 938 59200 994 60000 0 FreeSans 280 90 0 0 scan_in
port 5 nsew
flabel metal2 s 2870 59200 2926 60000 0 FreeSans 280 90 0 0 scan_out[0]
port 6 nsew
flabel metal2 s 22190 59200 22246 60000 0 FreeSans 280 90 0 0 scan_out[10]
port 7 nsew
flabel metal2 s 24122 59200 24178 60000 0 FreeSans 280 90 0 0 scan_out[11]
port 8 nsew
flabel metal2 s 26054 59200 26110 60000 0 FreeSans 280 90 0 0 scan_out[12]
port 9 nsew
flabel metal2 s 27986 59200 28042 60000 0 FreeSans 280 90 0 0 scan_out[13]
port 10 nsew
flabel metal2 s 29918 59200 29974 60000 0 FreeSans 280 90 0 0 scan_out[14]
port 11 nsew
flabel metal2 s 31850 59200 31906 60000 0 FreeSans 280 90 0 0 scan_out[15]
port 12 nsew
flabel metal2 s 33782 59200 33838 60000 0 FreeSans 280 90 0 0 scan_out[16]
port 13 nsew
flabel metal2 s 35714 59200 35770 60000 0 FreeSans 280 90 0 0 scan_out[17]
port 14 nsew
flabel metal2 s 37646 59200 37702 60000 0 FreeSans 280 90 0 0 scan_out[18]
port 15 nsew
flabel metal2 s 39578 59200 39634 60000 0 FreeSans 280 90 0 0 scan_out[19]
port 16 nsew
flabel metal2 s 4802 59200 4858 60000 0 FreeSans 280 90 0 0 scan_out[1]
port 17 nsew
flabel metal2 s 41510 59200 41566 60000 0 FreeSans 280 90 0 0 scan_out[20]
port 18 nsew
flabel metal2 s 43442 59200 43498 60000 0 FreeSans 280 90 0 0 scan_out[21]
port 19 nsew
flabel metal2 s 45374 59200 45430 60000 0 FreeSans 280 90 0 0 scan_out[22]
port 20 nsew
flabel metal2 s 47306 59200 47362 60000 0 FreeSans 280 90 0 0 scan_out[23]
port 21 nsew
flabel metal2 s 49238 59200 49294 60000 0 FreeSans 280 90 0 0 scan_out[24]
port 22 nsew
flabel metal2 s 51170 59200 51226 60000 0 FreeSans 280 90 0 0 scan_out[25]
port 23 nsew
flabel metal2 s 53102 59200 53158 60000 0 FreeSans 280 90 0 0 scan_out[26]
port 24 nsew
flabel metal2 s 55034 59200 55090 60000 0 FreeSans 280 90 0 0 scan_out[27]
port 25 nsew
flabel metal2 s 56966 59200 57022 60000 0 FreeSans 280 90 0 0 scan_out[28]
port 26 nsew
flabel metal2 s 58898 59200 58954 60000 0 FreeSans 280 90 0 0 scan_out[29]
port 27 nsew
flabel metal2 s 6734 59200 6790 60000 0 FreeSans 280 90 0 0 scan_out[2]
port 28 nsew
flabel metal2 s 8666 59200 8722 60000 0 FreeSans 280 90 0 0 scan_out[3]
port 29 nsew
flabel metal2 s 10598 59200 10654 60000 0 FreeSans 280 90 0 0 scan_out[4]
port 30 nsew
flabel metal2 s 12530 59200 12586 60000 0 FreeSans 280 90 0 0 scan_out[5]
port 31 nsew
flabel metal2 s 14462 59200 14518 60000 0 FreeSans 280 90 0 0 scan_out[6]
port 32 nsew
flabel metal2 s 16394 59200 16450 60000 0 FreeSans 280 90 0 0 scan_out[7]
port 33 nsew
flabel metal2 s 18326 59200 18382 60000 0 FreeSans 280 90 0 0 scan_out[8]
port 34 nsew
flabel metal2 s 20258 59200 20314 60000 0 FreeSans 280 90 0 0 scan_out[9]
port 35 nsew
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
