* NGSPICE file created from scan_chain.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

.subckt scan_chain VGND VPWR clk reset scan_in scan_out[0] scan_out[10] scan_out[11]
+ scan_out[12] scan_out[13] scan_out[14] scan_out[15] scan_out[16] scan_out[17] scan_out[18]
+ scan_out[19] scan_out[1] scan_out[20] scan_out[21] scan_out[22] scan_out[23] scan_out[24]
+ scan_out[25] scan_out[26] scan_out[27] scan_out[28] scan_out[29] scan_out[2] scan_out[3]
+ scan_out[4] scan_out[5] scan_out[6] scan_out[7] scan_out[8] scan_out[9]
XFILLER_0_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_131_ clknet_2_2__leaf_clk _005_ net43 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_114_ net4 net35 _032_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput20 net20 VGND VGND VPWR VPWR scan_out[25] sky130_fd_sc_hd__clkbuf_4
Xoutput7 net7 VGND VGND VPWR VPWR scan_out[13] sky130_fd_sc_hd__clkbuf_4
Xoutput31 net31 VGND VGND VPWR VPWR scan_out[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_130_ clknet_2_2__leaf_clk _004_ net43 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_113_ _036_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput21 net21 VGND VGND VPWR VPWR scan_out[26] sky130_fd_sc_hd__clkbuf_4
Xoutput10 net10 VGND VGND VPWR VPWR scan_out[16] sky130_fd_sc_hd__clkbuf_4
Xoutput8 net8 VGND VGND VPWR VPWR scan_out[14] sky130_fd_sc_hd__clkbuf_4
Xoutput32 net32 VGND VGND VPWR VPWR scan_out[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_112_ net32 net31 _032_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput22 net22 VGND VGND VPWR VPWR scan_out[27] sky130_fd_sc_hd__clkbuf_4
Xoutput11 net11 VGND VGND VPWR VPWR scan_out[17] sky130_fd_sc_hd__clkbuf_4
Xoutput9 net9 VGND VGND VPWR VPWR scan_out[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_111_ _035_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput23 net23 VGND VGND VPWR VPWR scan_out[28] sky130_fd_sc_hd__clkbuf_4
Xoutput12 net12 VGND VGND VPWR VPWR scan_out[18] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_110_ net31 net30 _032_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput24 net24 VGND VGND VPWR VPWR scan_out[29] sky130_fd_sc_hd__clkbuf_4
Xoutput13 net13 VGND VGND VPWR VPWR scan_out[19] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput25 net25 VGND VGND VPWR VPWR scan_out[2] sky130_fd_sc_hd__clkbuf_4
Xoutput14 net14 VGND VGND VPWR VPWR scan_out[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_099_ net26 net25 _053_ VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput15 net15 VGND VGND VPWR VPWR scan_out[20] sky130_fd_sc_hd__clkbuf_4
Xoutput26 net26 VGND VGND VPWR VPWR scan_out[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_098_ _061_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput16 net16 VGND VGND VPWR VPWR scan_out[21] sky130_fd_sc_hd__clkbuf_4
Xoutput27 net27 VGND VGND VPWR VPWR scan_out[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_84_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_097_ net25 net14 _053_ VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_149_ clknet_2_0__leaf_clk _023_ net41 VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput17 net17 VGND VGND VPWR VPWR scan_out[22] sky130_fd_sc_hd__clkbuf_4
Xoutput28 net28 VGND VGND VPWR VPWR scan_out[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_096_ _060_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_148_ clknet_2_0__leaf_clk _022_ net42 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_079_ _051_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput18 net18 VGND VGND VPWR VPWR scan_out[23] sky130_fd_sc_hd__clkbuf_4
Xoutput29 net29 VGND VGND VPWR VPWR scan_out[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_095_ net14 net3 _053_ VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_147_ clknet_2_1__leaf_clk _021_ net41 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_078_ net18 net34 _043_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput19 net19 VGND VGND VPWR VPWR scan_out[24] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_094_ _059_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_146_ clknet_2_0__leaf_clk _020_ net41 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_077_ _050_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_129_ clknet_2_2__leaf_clk _003_ net43 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_093_ _043_ net3 VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput1 reset VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_4
XFILLER_0_93_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_145_ clknet_2_1__leaf_clk _019_ net41 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dfrtp_1
X_076_ net34 net39 _043_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_128_ clknet_2_2__leaf_clk _002_ net43 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_092_ _058_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput2 scan_in VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_144_ clknet_2_0__leaf_clk _018_ net41 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_075_ _049_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_127_ clknet_2_1__leaf_clk _001_ net42 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_091_ net36 net23 _053_ VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_143_ clknet_2_0__leaf_clk _017_ net41 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_074_ net16 net15 _043_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_126_ clknet_2_1__leaf_clk _000_ net42 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_109_ _034_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_090_ _057_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_142_ clknet_2_1__leaf_clk _016_ net41 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_073_ _048_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_125_ _042_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_108_ net30 net29 _032_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_141_ clknet_2_1__leaf_clk _015_ net41 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_072_ net15 net13 _043_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_124_ net9 net33 _032_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_107_ _033_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_140_ clknet_2_0__leaf_clk _014_ net41 VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_071_ _047_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_123_ _041_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_106_ net29 net28 _032_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_070_ net13 net12 _043_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_122_ net8 net7 _032_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_105_ net2 VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_121_ net38 VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_104_ _031_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_120_ net7 net37 _032_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_103_ net28 net27 _053_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 net8 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_9_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_66_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_102_ _030_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2 net17 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_101_ net27 net26 _053_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 net32 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_100_ _062_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 net24 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold5 net6 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_089_ net23 net22 _053_ VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold6 _040_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_088_ _056_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold7 net16 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_087_ net22 net21 _053_ VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold8 net4 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_139_ clknet_2_3__leaf_clk _013_ net1 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_89_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_155_ clknet_2_1__leaf_clk _029_ net42 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_086_ _055_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_138_ clknet_2_3__leaf_clk _012_ net1 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_069_ _046_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_154_ clknet_2_0__leaf_clk _028_ net42 VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dfrtp_1
X_085_ net21 net20 _053_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_137_ clknet_2_3__leaf_clk _011_ net43 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_068_ net12 net11 _043_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout1 net42 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_153_ clknet_2_0__leaf_clk _027_ net42 VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_084_ _054_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_136_ clknet_2_3__leaf_clk _010_ net43 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_067_ _045_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_119_ _039_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout2 net1 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_152_ clknet_2_1__leaf_clk _026_ net42 VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_083_ net20 net19 _053_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_135_ clknet_2_3__leaf_clk _009_ net43 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_066_ net11 net10 _043_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_118_ net6 net5 _032_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout3 net1 VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput3 net3 VGND VGND VPWR VPWR scan_out[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_151_ clknet_2_1__leaf_clk _025_ net42 VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_082_ net2 VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__buf_4
XFILLER_0_33_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_134_ clknet_2_3__leaf_clk _008_ net43 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_065_ _044_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_117_ _038_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput4 net4 VGND VGND VPWR VPWR scan_out[10] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_150_ clknet_2_1__leaf_clk _024_ net41 VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_081_ _052_ VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_133_ clknet_2_3__leaf_clk _007_ net43 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_064_ net10 net9 _043_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_116_ net5 net40 _032_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput5 net5 VGND VGND VPWR VPWR scan_out[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_080_ net19 net18 _043_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_132_ clknet_2_2__leaf_clk _006_ net43 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_063_ net2 VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__buf_4
XFILLER_0_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_115_ _037_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput6 net6 VGND VGND VPWR VPWR scan_out[12] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput30 net30 VGND VGND VPWR VPWR scan_out[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
.ends

